VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO WB_InterConnect
  CLASS BLOCK ;
  FOREIGN WB_InterConnect ;
  ORIGIN 0.000 0.000 ;
  SIZE 1100.000 BY 1100.000 ;
  PIN clock
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.230 0.000 27.510 4.000 ;
    END
  END clock
  PIN io_dbus_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.760 4.000 20.360 ;
    END
  END io_dbus_addr[0]
  PIN io_dbus_addr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 223.760 4.000 224.360 ;
    END
  END io_dbus_addr[10]
  PIN io_dbus_addr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 240.760 4.000 241.360 ;
    END
  END io_dbus_addr[11]
  PIN io_dbus_addr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 258.440 4.000 259.040 ;
    END
  END io_dbus_addr[12]
  PIN io_dbus_addr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 276.120 4.000 276.720 ;
    END
  END io_dbus_addr[13]
  PIN io_dbus_addr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 293.800 4.000 294.400 ;
    END
  END io_dbus_addr[14]
  PIN io_dbus_addr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 310.800 4.000 311.400 ;
    END
  END io_dbus_addr[15]
  PIN io_dbus_addr[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 328.480 4.000 329.080 ;
    END
  END io_dbus_addr[16]
  PIN io_dbus_addr[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 346.160 4.000 346.760 ;
    END
  END io_dbus_addr[17]
  PIN io_dbus_addr[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 363.160 4.000 363.760 ;
    END
  END io_dbus_addr[18]
  PIN io_dbus_addr[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 380.840 4.000 381.440 ;
    END
  END io_dbus_addr[19]
  PIN io_dbus_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.000 4.000 49.600 ;
    END
  END io_dbus_addr[1]
  PIN io_dbus_addr[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 398.520 4.000 399.120 ;
    END
  END io_dbus_addr[20]
  PIN io_dbus_addr[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 415.520 4.000 416.120 ;
    END
  END io_dbus_addr[21]
  PIN io_dbus_addr[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 433.200 4.000 433.800 ;
    END
  END io_dbus_addr[22]
  PIN io_dbus_addr[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 450.880 4.000 451.480 ;
    END
  END io_dbus_addr[23]
  PIN io_dbus_addr[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 467.880 4.000 468.480 ;
    END
  END io_dbus_addr[24]
  PIN io_dbus_addr[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 485.560 4.000 486.160 ;
    END
  END io_dbus_addr[25]
  PIN io_dbus_addr[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 503.240 4.000 503.840 ;
    END
  END io_dbus_addr[26]
  PIN io_dbus_addr[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 520.240 4.000 520.840 ;
    END
  END io_dbus_addr[27]
  PIN io_dbus_addr[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 537.920 4.000 538.520 ;
    END
  END io_dbus_addr[28]
  PIN io_dbus_addr[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 555.600 4.000 556.200 ;
    END
  END io_dbus_addr[29]
  PIN io_dbus_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 4.000 78.840 ;
    END
  END io_dbus_addr[2]
  PIN io_dbus_addr[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 572.600 4.000 573.200 ;
    END
  END io_dbus_addr[30]
  PIN io_dbus_addr[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 590.280 4.000 590.880 ;
    END
  END io_dbus_addr[31]
  PIN io_dbus_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 101.360 4.000 101.960 ;
    END
  END io_dbus_addr[3]
  PIN io_dbus_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.040 4.000 119.640 ;
    END
  END io_dbus_addr[4]
  PIN io_dbus_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 4.000 136.640 ;
    END
  END io_dbus_addr[5]
  PIN io_dbus_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.720 4.000 154.320 ;
    END
  END io_dbus_addr[6]
  PIN io_dbus_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 171.400 4.000 172.000 ;
    END
  END io_dbus_addr[7]
  PIN io_dbus_addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 188.400 4.000 189.000 ;
    END
  END io_dbus_addr[8]
  PIN io_dbus_addr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 206.080 4.000 206.680 ;
    END
  END io_dbus_addr[9]
  PIN io_dbus_ld_type[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.880 4.000 26.480 ;
    END
  END io_dbus_ld_type[0]
  PIN io_dbus_ld_type[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.120 4.000 55.720 ;
    END
  END io_dbus_ld_type[1]
  PIN io_dbus_ld_type[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.680 4.000 84.280 ;
    END
  END io_dbus_ld_type[2]
  PIN io_dbus_rd_en
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.760 4.000 3.360 ;
    END
  END io_dbus_rd_en
  PIN io_dbus_rdata[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 31.320 4.000 31.920 ;
    END
  END io_dbus_rdata[0]
  PIN io_dbus_rdata[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 229.200 4.000 229.800 ;
    END
  END io_dbus_rdata[10]
  PIN io_dbus_rdata[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 246.880 4.000 247.480 ;
    END
  END io_dbus_rdata[11]
  PIN io_dbus_rdata[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 264.560 4.000 265.160 ;
    END
  END io_dbus_rdata[12]
  PIN io_dbus_rdata[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 281.560 4.000 282.160 ;
    END
  END io_dbus_rdata[13]
  PIN io_dbus_rdata[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 299.240 4.000 299.840 ;
    END
  END io_dbus_rdata[14]
  PIN io_dbus_rdata[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 316.920 4.000 317.520 ;
    END
  END io_dbus_rdata[15]
  PIN io_dbus_rdata[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 333.920 4.000 334.520 ;
    END
  END io_dbus_rdata[16]
  PIN io_dbus_rdata[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 351.600 4.000 352.200 ;
    END
  END io_dbus_rdata[17]
  PIN io_dbus_rdata[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 369.280 4.000 369.880 ;
    END
  END io_dbus_rdata[18]
  PIN io_dbus_rdata[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 386.960 4.000 387.560 ;
    END
  END io_dbus_rdata[19]
  PIN io_dbus_rdata[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 60.560 4.000 61.160 ;
    END
  END io_dbus_rdata[1]
  PIN io_dbus_rdata[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 403.960 4.000 404.560 ;
    END
  END io_dbus_rdata[20]
  PIN io_dbus_rdata[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 421.640 4.000 422.240 ;
    END
  END io_dbus_rdata[21]
  PIN io_dbus_rdata[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 439.320 4.000 439.920 ;
    END
  END io_dbus_rdata[22]
  PIN io_dbus_rdata[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 456.320 4.000 456.920 ;
    END
  END io_dbus_rdata[23]
  PIN io_dbus_rdata[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 474.000 4.000 474.600 ;
    END
  END io_dbus_rdata[24]
  PIN io_dbus_rdata[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 491.680 4.000 492.280 ;
    END
  END io_dbus_rdata[25]
  PIN io_dbus_rdata[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 508.680 4.000 509.280 ;
    END
  END io_dbus_rdata[26]
  PIN io_dbus_rdata[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 526.360 4.000 526.960 ;
    END
  END io_dbus_rdata[27]
  PIN io_dbus_rdata[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 544.040 4.000 544.640 ;
    END
  END io_dbus_rdata[28]
  PIN io_dbus_rdata[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 561.040 4.000 561.640 ;
    END
  END io_dbus_rdata[29]
  PIN io_dbus_rdata[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.800 4.000 90.400 ;
    END
  END io_dbus_rdata[2]
  PIN io_dbus_rdata[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 578.720 4.000 579.320 ;
    END
  END io_dbus_rdata[30]
  PIN io_dbus_rdata[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 596.400 4.000 597.000 ;
    END
  END io_dbus_rdata[31]
  PIN io_dbus_rdata[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 107.480 4.000 108.080 ;
    END
  END io_dbus_rdata[3]
  PIN io_dbus_rdata[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 124.480 4.000 125.080 ;
    END
  END io_dbus_rdata[4]
  PIN io_dbus_rdata[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.160 4.000 142.760 ;
    END
  END io_dbus_rdata[5]
  PIN io_dbus_rdata[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.840 4.000 160.440 ;
    END
  END io_dbus_rdata[6]
  PIN io_dbus_rdata[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.840 4.000 177.440 ;
    END
  END io_dbus_rdata[7]
  PIN io_dbus_rdata[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 194.520 4.000 195.120 ;
    END
  END io_dbus_rdata[8]
  PIN io_dbus_rdata[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 212.200 4.000 212.800 ;
    END
  END io_dbus_rdata[9]
  PIN io_dbus_st_type[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END io_dbus_st_type[0]
  PIN io_dbus_st_type[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.680 4.000 67.280 ;
    END
  END io_dbus_st_type[1]
  PIN io_dbus_valid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.200 4.000 8.800 ;
    END
  END io_dbus_valid
  PIN io_dbus_wdata[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.880 4.000 43.480 ;
    END
  END io_dbus_wdata[0]
  PIN io_dbus_wdata[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 235.320 4.000 235.920 ;
    END
  END io_dbus_wdata[10]
  PIN io_dbus_wdata[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 253.000 4.000 253.600 ;
    END
  END io_dbus_wdata[11]
  PIN io_dbus_wdata[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 270.000 4.000 270.600 ;
    END
  END io_dbus_wdata[12]
  PIN io_dbus_wdata[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 287.680 4.000 288.280 ;
    END
  END io_dbus_wdata[13]
  PIN io_dbus_wdata[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 305.360 4.000 305.960 ;
    END
  END io_dbus_wdata[14]
  PIN io_dbus_wdata[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 322.360 4.000 322.960 ;
    END
  END io_dbus_wdata[15]
  PIN io_dbus_wdata[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 340.040 4.000 340.640 ;
    END
  END io_dbus_wdata[16]
  PIN io_dbus_wdata[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 357.720 4.000 358.320 ;
    END
  END io_dbus_wdata[17]
  PIN io_dbus_wdata[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 374.720 4.000 375.320 ;
    END
  END io_dbus_wdata[18]
  PIN io_dbus_wdata[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 392.400 4.000 393.000 ;
    END
  END io_dbus_wdata[19]
  PIN io_dbus_wdata[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.120 4.000 72.720 ;
    END
  END io_dbus_wdata[1]
  PIN io_dbus_wdata[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 410.080 4.000 410.680 ;
    END
  END io_dbus_wdata[20]
  PIN io_dbus_wdata[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 427.080 4.000 427.680 ;
    END
  END io_dbus_wdata[21]
  PIN io_dbus_wdata[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 444.760 4.000 445.360 ;
    END
  END io_dbus_wdata[22]
  PIN io_dbus_wdata[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 462.440 4.000 463.040 ;
    END
  END io_dbus_wdata[23]
  PIN io_dbus_wdata[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 479.440 4.000 480.040 ;
    END
  END io_dbus_wdata[24]
  PIN io_dbus_wdata[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 497.120 4.000 497.720 ;
    END
  END io_dbus_wdata[25]
  PIN io_dbus_wdata[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 514.800 4.000 515.400 ;
    END
  END io_dbus_wdata[26]
  PIN io_dbus_wdata[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 532.480 4.000 533.080 ;
    END
  END io_dbus_wdata[27]
  PIN io_dbus_wdata[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 549.480 4.000 550.080 ;
    END
  END io_dbus_wdata[28]
  PIN io_dbus_wdata[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 567.160 4.000 567.760 ;
    END
  END io_dbus_wdata[29]
  PIN io_dbus_wdata[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END io_dbus_wdata[2]
  PIN io_dbus_wdata[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 584.840 4.000 585.440 ;
    END
  END io_dbus_wdata[30]
  PIN io_dbus_wdata[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 601.840 4.000 602.440 ;
    END
  END io_dbus_wdata[31]
  PIN io_dbus_wdata[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.920 4.000 113.520 ;
    END
  END io_dbus_wdata[3]
  PIN io_dbus_wdata[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 130.600 4.000 131.200 ;
    END
  END io_dbus_wdata[4]
  PIN io_dbus_wdata[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 148.280 4.000 148.880 ;
    END
  END io_dbus_wdata[5]
  PIN io_dbus_wdata[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 165.280 4.000 165.880 ;
    END
  END io_dbus_wdata[6]
  PIN io_dbus_wdata[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 182.960 4.000 183.560 ;
    END
  END io_dbus_wdata[7]
  PIN io_dbus_wdata[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 200.640 4.000 201.240 ;
    END
  END io_dbus_wdata[8]
  PIN io_dbus_wdata[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 217.640 4.000 218.240 ;
    END
  END io_dbus_wdata[9]
  PIN io_dbus_wr_en
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 14.320 4.000 14.920 ;
    END
  END io_dbus_wr_en
  PIN io_dmem_io_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.610 1096.000 28.890 1100.000 ;
    END
  END io_dmem_io_addr[0]
  PIN io_dmem_io_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.070 1096.000 75.350 1100.000 ;
    END
  END io_dmem_io_addr[1]
  PIN io_dmem_io_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.070 1096.000 121.350 1100.000 ;
    END
  END io_dmem_io_addr[2]
  PIN io_dmem_io_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 1096.000 167.810 1100.000 ;
    END
  END io_dmem_io_addr[3]
  PIN io_dmem_io_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.990 1096.000 214.270 1100.000 ;
    END
  END io_dmem_io_addr[4]
  PIN io_dmem_io_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.490 1096.000 248.770 1100.000 ;
    END
  END io_dmem_io_addr[5]
  PIN io_dmem_io_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.450 1096.000 283.730 1100.000 ;
    END
  END io_dmem_io_addr[6]
  PIN io_dmem_io_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.950 1096.000 318.230 1100.000 ;
    END
  END io_dmem_io_addr[7]
  PIN io_dmem_io_cs
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.610 1096.000 5.890 1100.000 ;
    END
  END io_dmem_io_cs
  PIN io_dmem_io_rdata[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.110 1096.000 40.390 1100.000 ;
    END
  END io_dmem_io_rdata[0]
  PIN io_dmem_io_rdata[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.910 1096.000 399.190 1100.000 ;
    END
  END io_dmem_io_rdata[10]
  PIN io_dmem_io_rdata[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 422.370 1096.000 422.650 1100.000 ;
    END
  END io_dmem_io_rdata[11]
  PIN io_dmem_io_rdata[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.370 1096.000 445.650 1100.000 ;
    END
  END io_dmem_io_rdata[12]
  PIN io_dmem_io_rdata[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 468.370 1096.000 468.650 1100.000 ;
    END
  END io_dmem_io_rdata[13]
  PIN io_dmem_io_rdata[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 491.830 1096.000 492.110 1100.000 ;
    END
  END io_dmem_io_rdata[14]
  PIN io_dmem_io_rdata[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 514.830 1096.000 515.110 1100.000 ;
    END
  END io_dmem_io_rdata[15]
  PIN io_dmem_io_rdata[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.830 1096.000 538.110 1100.000 ;
    END
  END io_dmem_io_rdata[16]
  PIN io_dmem_io_rdata[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 561.290 1096.000 561.570 1100.000 ;
    END
  END io_dmem_io_rdata[17]
  PIN io_dmem_io_rdata[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 584.290 1096.000 584.570 1100.000 ;
    END
  END io_dmem_io_rdata[18]
  PIN io_dmem_io_rdata[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 607.290 1096.000 607.570 1100.000 ;
    END
  END io_dmem_io_rdata[19]
  PIN io_dmem_io_rdata[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.570 1096.000 86.850 1100.000 ;
    END
  END io_dmem_io_rdata[1]
  PIN io_dmem_io_rdata[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 630.750 1096.000 631.030 1100.000 ;
    END
  END io_dmem_io_rdata[20]
  PIN io_dmem_io_rdata[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 653.750 1096.000 654.030 1100.000 ;
    END
  END io_dmem_io_rdata[21]
  PIN io_dmem_io_rdata[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 676.750 1096.000 677.030 1100.000 ;
    END
  END io_dmem_io_rdata[22]
  PIN io_dmem_io_rdata[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 700.210 1096.000 700.490 1100.000 ;
    END
  END io_dmem_io_rdata[23]
  PIN io_dmem_io_rdata[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 723.210 1096.000 723.490 1100.000 ;
    END
  END io_dmem_io_rdata[24]
  PIN io_dmem_io_rdata[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 746.210 1096.000 746.490 1100.000 ;
    END
  END io_dmem_io_rdata[25]
  PIN io_dmem_io_rdata[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 769.670 1096.000 769.950 1100.000 ;
    END
  END io_dmem_io_rdata[26]
  PIN io_dmem_io_rdata[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 792.670 1096.000 792.950 1100.000 ;
    END
  END io_dmem_io_rdata[27]
  PIN io_dmem_io_rdata[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 815.670 1096.000 815.950 1100.000 ;
    END
  END io_dmem_io_rdata[28]
  PIN io_dmem_io_rdata[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 839.130 1096.000 839.410 1100.000 ;
    END
  END io_dmem_io_rdata[29]
  PIN io_dmem_io_rdata[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.570 1096.000 132.850 1100.000 ;
    END
  END io_dmem_io_rdata[2]
  PIN io_dmem_io_rdata[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 862.130 1096.000 862.410 1100.000 ;
    END
  END io_dmem_io_rdata[30]
  PIN io_dmem_io_rdata[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 885.130 1096.000 885.410 1100.000 ;
    END
  END io_dmem_io_rdata[31]
  PIN io_dmem_io_rdata[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.030 1096.000 179.310 1100.000 ;
    END
  END io_dmem_io_rdata[3]
  PIN io_dmem_io_rdata[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.490 1096.000 225.770 1100.000 ;
    END
  END io_dmem_io_rdata[4]
  PIN io_dmem_io_rdata[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.990 1096.000 260.270 1100.000 ;
    END
  END io_dmem_io_rdata[5]
  PIN io_dmem_io_rdata[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.950 1096.000 295.230 1100.000 ;
    END
  END io_dmem_io_rdata[6]
  PIN io_dmem_io_rdata[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.450 1096.000 329.730 1100.000 ;
    END
  END io_dmem_io_rdata[7]
  PIN io_dmem_io_rdata[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 352.910 1096.000 353.190 1100.000 ;
    END
  END io_dmem_io_rdata[8]
  PIN io_dmem_io_rdata[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 375.910 1096.000 376.190 1100.000 ;
    END
  END io_dmem_io_rdata[9]
  PIN io_dmem_io_st_type[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 1096.000 51.890 1100.000 ;
    END
  END io_dmem_io_st_type[0]
  PIN io_dmem_io_st_type[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.070 1096.000 98.350 1100.000 ;
    END
  END io_dmem_io_st_type[1]
  PIN io_dmem_io_st_type[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.530 1096.000 144.810 1100.000 ;
    END
  END io_dmem_io_st_type[2]
  PIN io_dmem_io_st_type[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.530 1096.000 190.810 1100.000 ;
    END
  END io_dmem_io_st_type[3]
  PIN io_dmem_io_wdata[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.110 1096.000 63.390 1100.000 ;
    END
  END io_dmem_io_wdata[0]
  PIN io_dmem_io_wdata[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 410.410 1096.000 410.690 1100.000 ;
    END
  END io_dmem_io_wdata[10]
  PIN io_dmem_io_wdata[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 433.870 1096.000 434.150 1100.000 ;
    END
  END io_dmem_io_wdata[11]
  PIN io_dmem_io_wdata[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 456.870 1096.000 457.150 1100.000 ;
    END
  END io_dmem_io_wdata[12]
  PIN io_dmem_io_wdata[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.870 1096.000 480.150 1100.000 ;
    END
  END io_dmem_io_wdata[13]
  PIN io_dmem_io_wdata[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 503.330 1096.000 503.610 1100.000 ;
    END
  END io_dmem_io_wdata[14]
  PIN io_dmem_io_wdata[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 526.330 1096.000 526.610 1100.000 ;
    END
  END io_dmem_io_wdata[15]
  PIN io_dmem_io_wdata[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 549.330 1096.000 549.610 1100.000 ;
    END
  END io_dmem_io_wdata[16]
  PIN io_dmem_io_wdata[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 572.790 1096.000 573.070 1100.000 ;
    END
  END io_dmem_io_wdata[17]
  PIN io_dmem_io_wdata[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 595.790 1096.000 596.070 1100.000 ;
    END
  END io_dmem_io_wdata[18]
  PIN io_dmem_io_wdata[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 618.790 1096.000 619.070 1100.000 ;
    END
  END io_dmem_io_wdata[19]
  PIN io_dmem_io_wdata[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 1096.000 109.850 1100.000 ;
    END
  END io_dmem_io_wdata[1]
  PIN io_dmem_io_wdata[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 642.250 1096.000 642.530 1100.000 ;
    END
  END io_dmem_io_wdata[20]
  PIN io_dmem_io_wdata[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 665.250 1096.000 665.530 1100.000 ;
    END
  END io_dmem_io_wdata[21]
  PIN io_dmem_io_wdata[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 688.250 1096.000 688.530 1100.000 ;
    END
  END io_dmem_io_wdata[22]
  PIN io_dmem_io_wdata[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 711.710 1096.000 711.990 1100.000 ;
    END
  END io_dmem_io_wdata[23]
  PIN io_dmem_io_wdata[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 734.710 1096.000 734.990 1100.000 ;
    END
  END io_dmem_io_wdata[24]
  PIN io_dmem_io_wdata[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 757.710 1096.000 757.990 1100.000 ;
    END
  END io_dmem_io_wdata[25]
  PIN io_dmem_io_wdata[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 781.170 1096.000 781.450 1100.000 ;
    END
  END io_dmem_io_wdata[26]
  PIN io_dmem_io_wdata[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 804.170 1096.000 804.450 1100.000 ;
    END
  END io_dmem_io_wdata[27]
  PIN io_dmem_io_wdata[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 827.170 1096.000 827.450 1100.000 ;
    END
  END io_dmem_io_wdata[28]
  PIN io_dmem_io_wdata[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 850.630 1096.000 850.910 1100.000 ;
    END
  END io_dmem_io_wdata[29]
  PIN io_dmem_io_wdata[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.030 1096.000 156.310 1100.000 ;
    END
  END io_dmem_io_wdata[2]
  PIN io_dmem_io_wdata[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 873.630 1096.000 873.910 1100.000 ;
    END
  END io_dmem_io_wdata[30]
  PIN io_dmem_io_wdata[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 896.630 1096.000 896.910 1100.000 ;
    END
  END io_dmem_io_wdata[31]
  PIN io_dmem_io_wdata[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.030 1096.000 202.310 1100.000 ;
    END
  END io_dmem_io_wdata[3]
  PIN io_dmem_io_wdata[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.990 1096.000 237.270 1100.000 ;
    END
  END io_dmem_io_wdata[4]
  PIN io_dmem_io_wdata[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.490 1096.000 271.770 1100.000 ;
    END
  END io_dmem_io_wdata[5]
  PIN io_dmem_io_wdata[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 306.450 1096.000 306.730 1100.000 ;
    END
  END io_dmem_io_wdata[6]
  PIN io_dmem_io_wdata[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.950 1096.000 341.230 1100.000 ;
    END
  END io_dmem_io_wdata[7]
  PIN io_dmem_io_wdata[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 364.410 1096.000 364.690 1100.000 ;
    END
  END io_dmem_io_wdata[8]
  PIN io_dmem_io_wdata[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 387.410 1096.000 387.690 1100.000 ;
    END
  END io_dmem_io_wdata[9]
  PIN io_dmem_io_wr_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.110 1096.000 17.390 1100.000 ;
    END
  END io_dmem_io_wr_en
  PIN io_ibus_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 613.400 4.000 614.000 ;
    END
  END io_ibus_addr[0]
  PIN io_ibus_addr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 730.360 4.000 730.960 ;
    END
  END io_ibus_addr[10]
  PIN io_ibus_addr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 741.920 4.000 742.520 ;
    END
  END io_ibus_addr[11]
  PIN io_ibus_addr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 753.480 4.000 754.080 ;
    END
  END io_ibus_addr[12]
  PIN io_ibus_addr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 765.040 4.000 765.640 ;
    END
  END io_ibus_addr[13]
  PIN io_ibus_addr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 776.600 4.000 777.200 ;
    END
  END io_ibus_addr[14]
  PIN io_ibus_addr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 788.160 4.000 788.760 ;
    END
  END io_ibus_addr[15]
  PIN io_ibus_addr[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 799.720 4.000 800.320 ;
    END
  END io_ibus_addr[16]
  PIN io_ibus_addr[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 811.280 4.000 811.880 ;
    END
  END io_ibus_addr[17]
  PIN io_ibus_addr[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 823.520 4.000 824.120 ;
    END
  END io_ibus_addr[18]
  PIN io_ibus_addr[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 835.080 4.000 835.680 ;
    END
  END io_ibus_addr[19]
  PIN io_ibus_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 625.640 4.000 626.240 ;
    END
  END io_ibus_addr[1]
  PIN io_ibus_addr[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 846.640 4.000 847.240 ;
    END
  END io_ibus_addr[20]
  PIN io_ibus_addr[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 858.200 4.000 858.800 ;
    END
  END io_ibus_addr[21]
  PIN io_ibus_addr[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 869.760 4.000 870.360 ;
    END
  END io_ibus_addr[22]
  PIN io_ibus_addr[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 881.320 4.000 881.920 ;
    END
  END io_ibus_addr[23]
  PIN io_ibus_addr[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 892.880 4.000 893.480 ;
    END
  END io_ibus_addr[24]
  PIN io_ibus_addr[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 904.440 4.000 905.040 ;
    END
  END io_ibus_addr[25]
  PIN io_ibus_addr[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 916.680 4.000 917.280 ;
    END
  END io_ibus_addr[26]
  PIN io_ibus_addr[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 928.240 4.000 928.840 ;
    END
  END io_ibus_addr[27]
  PIN io_ibus_addr[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 939.800 4.000 940.400 ;
    END
  END io_ibus_addr[28]
  PIN io_ibus_addr[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 951.360 4.000 951.960 ;
    END
  END io_ibus_addr[29]
  PIN io_ibus_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 637.200 4.000 637.800 ;
    END
  END io_ibus_addr[2]
  PIN io_ibus_addr[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 962.920 4.000 963.520 ;
    END
  END io_ibus_addr[30]
  PIN io_ibus_addr[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 974.480 4.000 975.080 ;
    END
  END io_ibus_addr[31]
  PIN io_ibus_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 648.760 4.000 649.360 ;
    END
  END io_ibus_addr[3]
  PIN io_ibus_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 660.320 4.000 660.920 ;
    END
  END io_ibus_addr[4]
  PIN io_ibus_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 671.880 4.000 672.480 ;
    END
  END io_ibus_addr[5]
  PIN io_ibus_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 683.440 4.000 684.040 ;
    END
  END io_ibus_addr[6]
  PIN io_ibus_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 695.000 4.000 695.600 ;
    END
  END io_ibus_addr[7]
  PIN io_ibus_addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 706.560 4.000 707.160 ;
    END
  END io_ibus_addr[8]
  PIN io_ibus_addr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 718.120 4.000 718.720 ;
    END
  END io_ibus_addr[9]
  PIN io_ibus_inst[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 619.520 4.000 620.120 ;
    END
  END io_ibus_inst[0]
  PIN io_ibus_inst[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 735.800 4.000 736.400 ;
    END
  END io_ibus_inst[10]
  PIN io_ibus_inst[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 747.360 4.000 747.960 ;
    END
  END io_ibus_inst[11]
  PIN io_ibus_inst[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 758.920 4.000 759.520 ;
    END
  END io_ibus_inst[12]
  PIN io_ibus_inst[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 771.160 4.000 771.760 ;
    END
  END io_ibus_inst[13]
  PIN io_ibus_inst[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 782.720 4.000 783.320 ;
    END
  END io_ibus_inst[14]
  PIN io_ibus_inst[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 794.280 4.000 794.880 ;
    END
  END io_ibus_inst[15]
  PIN io_ibus_inst[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 805.840 4.000 806.440 ;
    END
  END io_ibus_inst[16]
  PIN io_ibus_inst[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 817.400 4.000 818.000 ;
    END
  END io_ibus_inst[17]
  PIN io_ibus_inst[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 828.960 4.000 829.560 ;
    END
  END io_ibus_inst[18]
  PIN io_ibus_inst[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 840.520 4.000 841.120 ;
    END
  END io_ibus_inst[19]
  PIN io_ibus_inst[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 631.080 4.000 631.680 ;
    END
  END io_ibus_inst[1]
  PIN io_ibus_inst[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 852.080 4.000 852.680 ;
    END
  END io_ibus_inst[20]
  PIN io_ibus_inst[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 864.320 4.000 864.920 ;
    END
  END io_ibus_inst[21]
  PIN io_ibus_inst[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 875.880 4.000 876.480 ;
    END
  END io_ibus_inst[22]
  PIN io_ibus_inst[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 887.440 4.000 888.040 ;
    END
  END io_ibus_inst[23]
  PIN io_ibus_inst[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 899.000 4.000 899.600 ;
    END
  END io_ibus_inst[24]
  PIN io_ibus_inst[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 910.560 4.000 911.160 ;
    END
  END io_ibus_inst[25]
  PIN io_ibus_inst[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 922.120 4.000 922.720 ;
    END
  END io_ibus_inst[26]
  PIN io_ibus_inst[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 933.680 4.000 934.280 ;
    END
  END io_ibus_inst[27]
  PIN io_ibus_inst[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 945.240 4.000 945.840 ;
    END
  END io_ibus_inst[28]
  PIN io_ibus_inst[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 956.800 4.000 957.400 ;
    END
  END io_ibus_inst[29]
  PIN io_ibus_inst[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 642.640 4.000 643.240 ;
    END
  END io_ibus_inst[2]
  PIN io_ibus_inst[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 969.040 4.000 969.640 ;
    END
  END io_ibus_inst[30]
  PIN io_ibus_inst[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 980.600 4.000 981.200 ;
    END
  END io_ibus_inst[31]
  PIN io_ibus_inst[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 654.200 4.000 654.800 ;
    END
  END io_ibus_inst[3]
  PIN io_ibus_inst[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 665.760 4.000 666.360 ;
    END
  END io_ibus_inst[4]
  PIN io_ibus_inst[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 678.000 4.000 678.600 ;
    END
  END io_ibus_inst[5]
  PIN io_ibus_inst[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 689.560 4.000 690.160 ;
    END
  END io_ibus_inst[6]
  PIN io_ibus_inst[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 701.120 4.000 701.720 ;
    END
  END io_ibus_inst[7]
  PIN io_ibus_inst[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 712.680 4.000 713.280 ;
    END
  END io_ibus_inst[8]
  PIN io_ibus_inst[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 724.240 4.000 724.840 ;
    END
  END io_ibus_inst[9]
  PIN io_ibus_valid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 607.960 4.000 608.560 ;
    END
  END io_ibus_valid
  PIN io_imem_io_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 876.560 1100.000 877.160 ;
    END
  END io_imem_io_addr[0]
  PIN io_imem_io_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.050 0.000 357.330 4.000 ;
    END
  END io_imem_io_addr[1]
  PIN io_imem_io_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 920.090 1096.000 920.370 1100.000 ;
    END
  END io_imem_io_addr[2]
  PIN io_imem_io_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1009.840 4.000 1010.440 ;
    END
  END io_imem_io_addr[3]
  PIN io_imem_io_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 895.600 1100.000 896.200 ;
    END
  END io_imem_io_addr[4]
  PIN io_imem_io_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 914.640 1100.000 915.240 ;
    END
  END io_imem_io_addr[5]
  PIN io_imem_io_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 933.000 1100.000 933.600 ;
    END
  END io_imem_io_addr[6]
  PIN io_imem_io_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 521.730 0.000 522.010 4.000 ;
    END
  END io_imem_io_addr[7]
  PIN io_imem_io_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.930 0.000 577.210 4.000 ;
    END
  END io_imem_io_addr[8]
  PIN io_imem_io_cs
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 908.590 1096.000 908.870 1100.000 ;
    END
  END io_imem_io_cs
  PIN io_imem_io_rdata[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.850 0.000 302.130 4.000 ;
    END
  END io_imem_io_rdata[0]
  PIN io_imem_io_rdata[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 971.080 1100.000 971.680 ;
    END
  END io_imem_io_rdata[10]
  PIN io_imem_io_rdata[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 980.600 1100.000 981.200 ;
    END
  END io_imem_io_rdata[11]
  PIN io_imem_io_rdata[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 990.120 1100.000 990.720 ;
    END
  END io_imem_io_rdata[12]
  PIN io_imem_io_rdata[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1044.520 4.000 1045.120 ;
    END
  END io_imem_io_rdata[13]
  PIN io_imem_io_rdata[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1049.960 4.000 1050.560 ;
    END
  END io_imem_io_rdata[14]
  PIN io_imem_io_rdata[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 1009.160 1100.000 1009.760 ;
    END
  END io_imem_io_rdata[15]
  PIN io_imem_io_rdata[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 686.870 0.000 687.150 4.000 ;
    END
  END io_imem_io_rdata[16]
  PIN io_imem_io_rdata[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 1018.680 1100.000 1019.280 ;
    END
  END io_imem_io_rdata[17]
  PIN io_imem_io_rdata[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1062.200 4.000 1062.800 ;
    END
  END io_imem_io_rdata[18]
  PIN io_imem_io_rdata[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1067.640 4.000 1068.240 ;
    END
  END io_imem_io_rdata[19]
  PIN io_imem_io_rdata[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 411.790 0.000 412.070 4.000 ;
    END
  END io_imem_io_rdata[1]
  PIN io_imem_io_rdata[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1073.760 4.000 1074.360 ;
    END
  END io_imem_io_rdata[20]
  PIN io_imem_io_rdata[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1024.050 1096.000 1024.330 1100.000 ;
    END
  END io_imem_io_rdata[21]
  PIN io_imem_io_rdata[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1085.320 4.000 1085.920 ;
    END
  END io_imem_io_rdata[22]
  PIN io_imem_io_rdata[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1090.760 4.000 1091.360 ;
    END
  END io_imem_io_rdata[23]
  PIN io_imem_io_rdata[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1035.550 1096.000 1035.830 1100.000 ;
    END
  END io_imem_io_rdata[24]
  PIN io_imem_io_rdata[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 961.950 0.000 962.230 4.000 ;
    END
  END io_imem_io_rdata[25]
  PIN io_imem_io_rdata[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 1056.760 1100.000 1057.360 ;
    END
  END io_imem_io_rdata[26]
  PIN io_imem_io_rdata[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1016.690 0.000 1016.970 4.000 ;
    END
  END io_imem_io_rdata[27]
  PIN io_imem_io_rdata[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1059.010 1096.000 1059.290 1100.000 ;
    END
  END io_imem_io_rdata[28]
  PIN io_imem_io_rdata[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1096.880 4.000 1097.480 ;
    END
  END io_imem_io_rdata[29]
  PIN io_imem_io_rdata[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 931.590 1096.000 931.870 1100.000 ;
    END
  END io_imem_io_rdata[2]
  PIN io_imem_io_rdata[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1070.510 1096.000 1070.790 1100.000 ;
    END
  END io_imem_io_rdata[30]
  PIN io_imem_io_rdata[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1071.890 0.000 1072.170 4.000 ;
    END
  END io_imem_io_rdata[31]
  PIN io_imem_io_rdata[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 886.080 1100.000 886.680 ;
    END
  END io_imem_io_rdata[3]
  PIN io_imem_io_rdata[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 905.120 1100.000 905.720 ;
    END
  END io_imem_io_rdata[4]
  PIN io_imem_io_rdata[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 923.480 1100.000 924.080 ;
    END
  END io_imem_io_rdata[5]
  PIN io_imem_io_rdata[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1015.280 4.000 1015.880 ;
    END
  END io_imem_io_rdata[6]
  PIN io_imem_io_rdata[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1021.400 4.000 1022.000 ;
    END
  END io_imem_io_rdata[7]
  PIN io_imem_io_rdata[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 989.550 1096.000 989.830 1100.000 ;
    END
  END io_imem_io_rdata[8]
  PIN io_imem_io_rdata[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1026.840 4.000 1027.440 ;
    END
  END io_imem_io_rdata[9]
  PIN io_imem_io_wdata[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 997.600 4.000 998.200 ;
    END
  END io_imem_io_wdata[0]
  PIN io_imem_io_wdata[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1032.960 4.000 1033.560 ;
    END
  END io_imem_io_wdata[10]
  PIN io_imem_io_wdata[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1001.050 1096.000 1001.330 1100.000 ;
    END
  END io_imem_io_wdata[11]
  PIN io_imem_io_wdata[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1038.400 4.000 1039.000 ;
    END
  END io_imem_io_wdata[12]
  PIN io_imem_io_wdata[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 999.640 1100.000 1000.240 ;
    END
  END io_imem_io_wdata[13]
  PIN io_imem_io_wdata[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1056.080 4.000 1056.680 ;
    END
  END io_imem_io_wdata[14]
  PIN io_imem_io_wdata[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 632.130 0.000 632.410 4.000 ;
    END
  END io_imem_io_wdata[15]
  PIN io_imem_io_wdata[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1012.550 1096.000 1012.830 1100.000 ;
    END
  END io_imem_io_wdata[16]
  PIN io_imem_io_wdata[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 742.070 0.000 742.350 4.000 ;
    END
  END io_imem_io_wdata[17]
  PIN io_imem_io_wdata[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 796.810 0.000 797.090 4.000 ;
    END
  END io_imem_io_wdata[18]
  PIN io_imem_io_wdata[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 852.010 0.000 852.290 4.000 ;
    END
  END io_imem_io_wdata[19]
  PIN io_imem_io_wdata[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1003.720 4.000 1004.320 ;
    END
  END io_imem_io_wdata[1]
  PIN io_imem_io_wdata[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1079.200 4.000 1079.800 ;
    END
  END io_imem_io_wdata[20]
  PIN io_imem_io_wdata[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 1028.200 1100.000 1028.800 ;
    END
  END io_imem_io_wdata[21]
  PIN io_imem_io_wdata[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 906.750 0.000 907.030 4.000 ;
    END
  END io_imem_io_wdata[22]
  PIN io_imem_io_wdata[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 1037.720 1100.000 1038.320 ;
    END
  END io_imem_io_wdata[23]
  PIN io_imem_io_wdata[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1047.510 1096.000 1047.790 1100.000 ;
    END
  END io_imem_io_wdata[24]
  PIN io_imem_io_wdata[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 1047.240 1100.000 1047.840 ;
    END
  END io_imem_io_wdata[25]
  PIN io_imem_io_wdata[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 1066.280 1100.000 1066.880 ;
    END
  END io_imem_io_wdata[26]
  PIN io_imem_io_wdata[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 1075.800 1100.000 1076.400 ;
    END
  END io_imem_io_wdata[27]
  PIN io_imem_io_wdata[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 1085.320 1100.000 1085.920 ;
    END
  END io_imem_io_wdata[28]
  PIN io_imem_io_wdata[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 1094.840 1100.000 1095.440 ;
    END
  END io_imem_io_wdata[29]
  PIN io_imem_io_wdata[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 943.090 1096.000 943.370 1100.000 ;
    END
  END io_imem_io_wdata[2]
  PIN io_imem_io_wdata[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1082.010 1096.000 1082.290 1100.000 ;
    END
  END io_imem_io_wdata[30]
  PIN io_imem_io_wdata[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1093.510 1096.000 1093.790 1100.000 ;
    END
  END io_imem_io_wdata[31]
  PIN io_imem_io_wdata[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.990 0.000 467.270 4.000 ;
    END
  END io_imem_io_wdata[3]
  PIN io_imem_io_wdata[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 954.590 1096.000 954.870 1100.000 ;
    END
  END io_imem_io_wdata[4]
  PIN io_imem_io_wdata[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 966.090 1096.000 966.370 1100.000 ;
    END
  END io_imem_io_wdata[5]
  PIN io_imem_io_wdata[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 942.520 1100.000 943.120 ;
    END
  END io_imem_io_wdata[6]
  PIN io_imem_io_wdata[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 978.050 1096.000 978.330 1100.000 ;
    END
  END io_imem_io_wdata[7]
  PIN io_imem_io_wdata[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 952.040 1100.000 952.640 ;
    END
  END io_imem_io_wdata[8]
  PIN io_imem_io_wdata[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 961.560 1100.000 962.160 ;
    END
  END io_imem_io_wdata[9]
  PIN io_imem_io_wr_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.110 0.000 247.390 4.000 ;
    END
  END io_imem_io_wr_en
  PIN io_motor_ack_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 4.120 1100.000 4.720 ;
    END
  END io_motor_ack_i
  PIN io_motor_addr_sel
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 12.960 1100.000 13.560 ;
    END
  END io_motor_addr_sel
  PIN io_motor_data_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 22.480 1100.000 23.080 ;
    END
  END io_motor_data_i[0]
  PIN io_motor_data_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 117.680 1100.000 118.280 ;
    END
  END io_motor_data_i[10]
  PIN io_motor_data_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 127.200 1100.000 127.800 ;
    END
  END io_motor_data_i[11]
  PIN io_motor_data_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 136.720 1100.000 137.320 ;
    END
  END io_motor_data_i[12]
  PIN io_motor_data_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 146.240 1100.000 146.840 ;
    END
  END io_motor_data_i[13]
  PIN io_motor_data_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 155.760 1100.000 156.360 ;
    END
  END io_motor_data_i[14]
  PIN io_motor_data_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 165.280 1100.000 165.880 ;
    END
  END io_motor_data_i[15]
  PIN io_motor_data_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 174.800 1100.000 175.400 ;
    END
  END io_motor_data_i[16]
  PIN io_motor_data_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 184.320 1100.000 184.920 ;
    END
  END io_motor_data_i[17]
  PIN io_motor_data_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 193.160 1100.000 193.760 ;
    END
  END io_motor_data_i[18]
  PIN io_motor_data_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 202.680 1100.000 203.280 ;
    END
  END io_motor_data_i[19]
  PIN io_motor_data_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 32.000 1100.000 32.600 ;
    END
  END io_motor_data_i[1]
  PIN io_motor_data_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 212.200 1100.000 212.800 ;
    END
  END io_motor_data_i[20]
  PIN io_motor_data_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 221.720 1100.000 222.320 ;
    END
  END io_motor_data_i[21]
  PIN io_motor_data_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 231.240 1100.000 231.840 ;
    END
  END io_motor_data_i[22]
  PIN io_motor_data_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 240.760 1100.000 241.360 ;
    END
  END io_motor_data_i[23]
  PIN io_motor_data_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 250.280 1100.000 250.880 ;
    END
  END io_motor_data_i[24]
  PIN io_motor_data_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 259.800 1100.000 260.400 ;
    END
  END io_motor_data_i[25]
  PIN io_motor_data_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 269.320 1100.000 269.920 ;
    END
  END io_motor_data_i[26]
  PIN io_motor_data_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 278.840 1100.000 279.440 ;
    END
  END io_motor_data_i[27]
  PIN io_motor_data_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 288.360 1100.000 288.960 ;
    END
  END io_motor_data_i[28]
  PIN io_motor_data_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 297.880 1100.000 298.480 ;
    END
  END io_motor_data_i[29]
  PIN io_motor_data_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 41.520 1100.000 42.120 ;
    END
  END io_motor_data_i[2]
  PIN io_motor_data_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 307.400 1100.000 308.000 ;
    END
  END io_motor_data_i[30]
  PIN io_motor_data_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 316.920 1100.000 317.520 ;
    END
  END io_motor_data_i[31]
  PIN io_motor_data_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 51.040 1100.000 51.640 ;
    END
  END io_motor_data_i[3]
  PIN io_motor_data_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 60.560 1100.000 61.160 ;
    END
  END io_motor_data_i[4]
  PIN io_motor_data_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 70.080 1100.000 70.680 ;
    END
  END io_motor_data_i[5]
  PIN io_motor_data_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 79.600 1100.000 80.200 ;
    END
  END io_motor_data_i[6]
  PIN io_motor_data_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 89.120 1100.000 89.720 ;
    END
  END io_motor_data_i[7]
  PIN io_motor_data_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 98.640 1100.000 99.240 ;
    END
  END io_motor_data_i[8]
  PIN io_motor_data_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 108.160 1100.000 108.760 ;
    END
  END io_motor_data_i[9]
  PIN io_spi_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 838.480 1100.000 839.080 ;
    END
  END io_spi_clk
  PIN io_spi_cs
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 848.000 1100.000 848.600 ;
    END
  END io_spi_cs
  PIN io_spi_irq
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 986.040 4.000 986.640 ;
    END
  END io_spi_irq
  PIN io_spi_miso
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.170 0.000 137.450 4.000 ;
    END
  END io_spi_miso
  PIN io_spi_mosi
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 857.520 1100.000 858.120 ;
    END
  END io_spi_mosi
  PIN io_uart_irq
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 992.160 4.000 992.760 ;
    END
  END io_uart_irq
  PIN io_uart_rx
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.910 0.000 192.190 4.000 ;
    END
  END io_uart_rx
  PIN io_uart_tx
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 867.040 1100.000 867.640 ;
    END
  END io_uart_tx
  PIN io_wbm_m2s_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 345.480 1100.000 346.080 ;
    END
  END io_wbm_m2s_addr[0]
  PIN io_wbm_m2s_addr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 572.600 1100.000 573.200 ;
    END
  END io_wbm_m2s_addr[10]
  PIN io_wbm_m2s_addr[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 591.640 1100.000 592.240 ;
    END
  END io_wbm_m2s_addr[11]
  PIN io_wbm_m2s_addr[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 610.680 1100.000 611.280 ;
    END
  END io_wbm_m2s_addr[12]
  PIN io_wbm_m2s_addr[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 629.720 1100.000 630.320 ;
    END
  END io_wbm_m2s_addr[13]
  PIN io_wbm_m2s_addr[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 648.760 1100.000 649.360 ;
    END
  END io_wbm_m2s_addr[14]
  PIN io_wbm_m2s_addr[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 667.800 1100.000 668.400 ;
    END
  END io_wbm_m2s_addr[15]
  PIN io_wbm_m2s_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 373.360 1100.000 373.960 ;
    END
  END io_wbm_m2s_addr[1]
  PIN io_wbm_m2s_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 401.920 1100.000 402.520 ;
    END
  END io_wbm_m2s_addr[2]
  PIN io_wbm_m2s_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 430.480 1100.000 431.080 ;
    END
  END io_wbm_m2s_addr[3]
  PIN io_wbm_m2s_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 459.040 1100.000 459.640 ;
    END
  END io_wbm_m2s_addr[4]
  PIN io_wbm_m2s_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 478.080 1100.000 478.680 ;
    END
  END io_wbm_m2s_addr[5]
  PIN io_wbm_m2s_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 497.120 1100.000 497.720 ;
    END
  END io_wbm_m2s_addr[6]
  PIN io_wbm_m2s_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 516.160 1100.000 516.760 ;
    END
  END io_wbm_m2s_addr[7]
  PIN io_wbm_m2s_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 535.200 1100.000 535.800 ;
    END
  END io_wbm_m2s_addr[8]
  PIN io_wbm_m2s_addr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 554.240 1100.000 554.840 ;
    END
  END io_wbm_m2s_addr[9]
  PIN io_wbm_m2s_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 355.000 1100.000 355.600 ;
    END
  END io_wbm_m2s_data[0]
  PIN io_wbm_m2s_data[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 582.120 1100.000 582.720 ;
    END
  END io_wbm_m2s_data[10]
  PIN io_wbm_m2s_data[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 601.160 1100.000 601.760 ;
    END
  END io_wbm_m2s_data[11]
  PIN io_wbm_m2s_data[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 620.200 1100.000 620.800 ;
    END
  END io_wbm_m2s_data[12]
  PIN io_wbm_m2s_data[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 639.240 1100.000 639.840 ;
    END
  END io_wbm_m2s_data[13]
  PIN io_wbm_m2s_data[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 658.280 1100.000 658.880 ;
    END
  END io_wbm_m2s_data[14]
  PIN io_wbm_m2s_data[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 677.320 1100.000 677.920 ;
    END
  END io_wbm_m2s_data[15]
  PIN io_wbm_m2s_data[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 686.840 1100.000 687.440 ;
    END
  END io_wbm_m2s_data[16]
  PIN io_wbm_m2s_data[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 696.360 1100.000 696.960 ;
    END
  END io_wbm_m2s_data[17]
  PIN io_wbm_m2s_data[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 705.880 1100.000 706.480 ;
    END
  END io_wbm_m2s_data[18]
  PIN io_wbm_m2s_data[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 715.400 1100.000 716.000 ;
    END
  END io_wbm_m2s_data[19]
  PIN io_wbm_m2s_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 382.880 1100.000 383.480 ;
    END
  END io_wbm_m2s_data[1]
  PIN io_wbm_m2s_data[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 724.920 1100.000 725.520 ;
    END
  END io_wbm_m2s_data[20]
  PIN io_wbm_m2s_data[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 734.440 1100.000 735.040 ;
    END
  END io_wbm_m2s_data[21]
  PIN io_wbm_m2s_data[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 743.280 1100.000 743.880 ;
    END
  END io_wbm_m2s_data[22]
  PIN io_wbm_m2s_data[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 752.800 1100.000 753.400 ;
    END
  END io_wbm_m2s_data[23]
  PIN io_wbm_m2s_data[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 762.320 1100.000 762.920 ;
    END
  END io_wbm_m2s_data[24]
  PIN io_wbm_m2s_data[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 771.840 1100.000 772.440 ;
    END
  END io_wbm_m2s_data[25]
  PIN io_wbm_m2s_data[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 781.360 1100.000 781.960 ;
    END
  END io_wbm_m2s_data[26]
  PIN io_wbm_m2s_data[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 790.880 1100.000 791.480 ;
    END
  END io_wbm_m2s_data[27]
  PIN io_wbm_m2s_data[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 800.400 1100.000 801.000 ;
    END
  END io_wbm_m2s_data[28]
  PIN io_wbm_m2s_data[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 809.920 1100.000 810.520 ;
    END
  END io_wbm_m2s_data[29]
  PIN io_wbm_m2s_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 411.440 1100.000 412.040 ;
    END
  END io_wbm_m2s_data[2]
  PIN io_wbm_m2s_data[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 819.440 1100.000 820.040 ;
    END
  END io_wbm_m2s_data[30]
  PIN io_wbm_m2s_data[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 828.960 1100.000 829.560 ;
    END
  END io_wbm_m2s_data[31]
  PIN io_wbm_m2s_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 440.000 1100.000 440.600 ;
    END
  END io_wbm_m2s_data[3]
  PIN io_wbm_m2s_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 468.560 1100.000 469.160 ;
    END
  END io_wbm_m2s_data[4]
  PIN io_wbm_m2s_data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 487.600 1100.000 488.200 ;
    END
  END io_wbm_m2s_data[5]
  PIN io_wbm_m2s_data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 506.640 1100.000 507.240 ;
    END
  END io_wbm_m2s_data[6]
  PIN io_wbm_m2s_data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 525.680 1100.000 526.280 ;
    END
  END io_wbm_m2s_data[7]
  PIN io_wbm_m2s_data[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 544.720 1100.000 545.320 ;
    END
  END io_wbm_m2s_data[8]
  PIN io_wbm_m2s_data[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 563.080 1100.000 563.680 ;
    END
  END io_wbm_m2s_data[9]
  PIN io_wbm_m2s_sel[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 364.520 1100.000 365.120 ;
    END
  END io_wbm_m2s_sel[0]
  PIN io_wbm_m2s_sel[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 392.400 1100.000 393.000 ;
    END
  END io_wbm_m2s_sel[1]
  PIN io_wbm_m2s_sel[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 420.960 1100.000 421.560 ;
    END
  END io_wbm_m2s_sel[2]
  PIN io_wbm_m2s_sel[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 449.520 1100.000 450.120 ;
    END
  END io_wbm_m2s_sel[3]
  PIN io_wbm_m2s_stb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 326.440 1100.000 327.040 ;
    END
  END io_wbm_m2s_stb
  PIN io_wbm_m2s_we
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 335.960 1100.000 336.560 ;
    END
  END io_wbm_m2s_we
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.970 0.000 82.250 4.000 ;
    END
  END reset
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1088.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 1088.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 1088.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 1088.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 1088.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 1088.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 1088.240 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1088.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 1088.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 1088.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 1088.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 1088.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 1088.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 1088.240 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 1094.340 1088.085 ;
      LAYER met1 ;
        RECT 5.520 10.640 1094.340 1088.980 ;
      LAYER met2 ;
        RECT 6.170 1095.720 16.830 1097.365 ;
        RECT 17.670 1095.720 28.330 1097.365 ;
        RECT 29.170 1095.720 39.830 1097.365 ;
        RECT 40.670 1095.720 51.330 1097.365 ;
        RECT 52.170 1095.720 62.830 1097.365 ;
        RECT 63.670 1095.720 74.790 1097.365 ;
        RECT 75.630 1095.720 86.290 1097.365 ;
        RECT 87.130 1095.720 97.790 1097.365 ;
        RECT 98.630 1095.720 109.290 1097.365 ;
        RECT 110.130 1095.720 120.790 1097.365 ;
        RECT 121.630 1095.720 132.290 1097.365 ;
        RECT 133.130 1095.720 144.250 1097.365 ;
        RECT 145.090 1095.720 155.750 1097.365 ;
        RECT 156.590 1095.720 167.250 1097.365 ;
        RECT 168.090 1095.720 178.750 1097.365 ;
        RECT 179.590 1095.720 190.250 1097.365 ;
        RECT 191.090 1095.720 201.750 1097.365 ;
        RECT 202.590 1095.720 213.710 1097.365 ;
        RECT 214.550 1095.720 225.210 1097.365 ;
        RECT 226.050 1095.720 236.710 1097.365 ;
        RECT 237.550 1095.720 248.210 1097.365 ;
        RECT 249.050 1095.720 259.710 1097.365 ;
        RECT 260.550 1095.720 271.210 1097.365 ;
        RECT 272.050 1095.720 283.170 1097.365 ;
        RECT 284.010 1095.720 294.670 1097.365 ;
        RECT 295.510 1095.720 306.170 1097.365 ;
        RECT 307.010 1095.720 317.670 1097.365 ;
        RECT 318.510 1095.720 329.170 1097.365 ;
        RECT 330.010 1095.720 340.670 1097.365 ;
        RECT 341.510 1095.720 352.630 1097.365 ;
        RECT 353.470 1095.720 364.130 1097.365 ;
        RECT 364.970 1095.720 375.630 1097.365 ;
        RECT 376.470 1095.720 387.130 1097.365 ;
        RECT 387.970 1095.720 398.630 1097.365 ;
        RECT 399.470 1095.720 410.130 1097.365 ;
        RECT 410.970 1095.720 422.090 1097.365 ;
        RECT 422.930 1095.720 433.590 1097.365 ;
        RECT 434.430 1095.720 445.090 1097.365 ;
        RECT 445.930 1095.720 456.590 1097.365 ;
        RECT 457.430 1095.720 468.090 1097.365 ;
        RECT 468.930 1095.720 479.590 1097.365 ;
        RECT 480.430 1095.720 491.550 1097.365 ;
        RECT 492.390 1095.720 503.050 1097.365 ;
        RECT 503.890 1095.720 514.550 1097.365 ;
        RECT 515.390 1095.720 526.050 1097.365 ;
        RECT 526.890 1095.720 537.550 1097.365 ;
        RECT 538.390 1095.720 549.050 1097.365 ;
        RECT 549.890 1095.720 561.010 1097.365 ;
        RECT 561.850 1095.720 572.510 1097.365 ;
        RECT 573.350 1095.720 584.010 1097.365 ;
        RECT 584.850 1095.720 595.510 1097.365 ;
        RECT 596.350 1095.720 607.010 1097.365 ;
        RECT 607.850 1095.720 618.510 1097.365 ;
        RECT 619.350 1095.720 630.470 1097.365 ;
        RECT 631.310 1095.720 641.970 1097.365 ;
        RECT 642.810 1095.720 653.470 1097.365 ;
        RECT 654.310 1095.720 664.970 1097.365 ;
        RECT 665.810 1095.720 676.470 1097.365 ;
        RECT 677.310 1095.720 687.970 1097.365 ;
        RECT 688.810 1095.720 699.930 1097.365 ;
        RECT 700.770 1095.720 711.430 1097.365 ;
        RECT 712.270 1095.720 722.930 1097.365 ;
        RECT 723.770 1095.720 734.430 1097.365 ;
        RECT 735.270 1095.720 745.930 1097.365 ;
        RECT 746.770 1095.720 757.430 1097.365 ;
        RECT 758.270 1095.720 769.390 1097.365 ;
        RECT 770.230 1095.720 780.890 1097.365 ;
        RECT 781.730 1095.720 792.390 1097.365 ;
        RECT 793.230 1095.720 803.890 1097.365 ;
        RECT 804.730 1095.720 815.390 1097.365 ;
        RECT 816.230 1095.720 826.890 1097.365 ;
        RECT 827.730 1095.720 838.850 1097.365 ;
        RECT 839.690 1095.720 850.350 1097.365 ;
        RECT 851.190 1095.720 861.850 1097.365 ;
        RECT 862.690 1095.720 873.350 1097.365 ;
        RECT 874.190 1095.720 884.850 1097.365 ;
        RECT 885.690 1095.720 896.350 1097.365 ;
        RECT 897.190 1095.720 908.310 1097.365 ;
        RECT 909.150 1095.720 919.810 1097.365 ;
        RECT 920.650 1095.720 931.310 1097.365 ;
        RECT 932.150 1095.720 942.810 1097.365 ;
        RECT 943.650 1095.720 954.310 1097.365 ;
        RECT 955.150 1095.720 965.810 1097.365 ;
        RECT 966.650 1095.720 977.770 1097.365 ;
        RECT 978.610 1095.720 989.270 1097.365 ;
        RECT 990.110 1095.720 1000.770 1097.365 ;
        RECT 1001.610 1095.720 1012.270 1097.365 ;
        RECT 1013.110 1095.720 1023.770 1097.365 ;
        RECT 1024.610 1095.720 1035.270 1097.365 ;
        RECT 1036.110 1095.720 1047.230 1097.365 ;
        RECT 1048.070 1095.720 1058.730 1097.365 ;
        RECT 1059.570 1095.720 1070.230 1097.365 ;
        RECT 1071.070 1095.720 1081.730 1097.365 ;
        RECT 1082.570 1095.720 1093.230 1097.365 ;
        RECT 5.620 4.280 1093.780 1095.720 ;
        RECT 5.620 2.875 26.950 4.280 ;
        RECT 27.790 2.875 81.690 4.280 ;
        RECT 82.530 2.875 136.890 4.280 ;
        RECT 137.730 2.875 191.630 4.280 ;
        RECT 192.470 2.875 246.830 4.280 ;
        RECT 247.670 2.875 301.570 4.280 ;
        RECT 302.410 2.875 356.770 4.280 ;
        RECT 357.610 2.875 411.510 4.280 ;
        RECT 412.350 2.875 466.710 4.280 ;
        RECT 467.550 2.875 521.450 4.280 ;
        RECT 522.290 2.875 576.650 4.280 ;
        RECT 577.490 2.875 631.850 4.280 ;
        RECT 632.690 2.875 686.590 4.280 ;
        RECT 687.430 2.875 741.790 4.280 ;
        RECT 742.630 2.875 796.530 4.280 ;
        RECT 797.370 2.875 851.730 4.280 ;
        RECT 852.570 2.875 906.470 4.280 ;
        RECT 907.310 2.875 961.670 4.280 ;
        RECT 962.510 2.875 1016.410 4.280 ;
        RECT 1017.250 2.875 1071.610 4.280 ;
        RECT 1072.450 2.875 1093.780 4.280 ;
      LAYER met3 ;
        RECT 4.400 1096.480 1096.000 1097.345 ;
        RECT 4.000 1095.840 1096.000 1096.480 ;
        RECT 4.000 1094.440 1095.600 1095.840 ;
        RECT 4.000 1091.760 1096.000 1094.440 ;
        RECT 4.400 1090.360 1096.000 1091.760 ;
        RECT 4.000 1086.320 1096.000 1090.360 ;
        RECT 4.400 1084.920 1095.600 1086.320 ;
        RECT 4.000 1080.200 1096.000 1084.920 ;
        RECT 4.400 1078.800 1096.000 1080.200 ;
        RECT 4.000 1076.800 1096.000 1078.800 ;
        RECT 4.000 1075.400 1095.600 1076.800 ;
        RECT 4.000 1074.760 1096.000 1075.400 ;
        RECT 4.400 1073.360 1096.000 1074.760 ;
        RECT 4.000 1068.640 1096.000 1073.360 ;
        RECT 4.400 1067.280 1096.000 1068.640 ;
        RECT 4.400 1067.240 1095.600 1067.280 ;
        RECT 4.000 1065.880 1095.600 1067.240 ;
        RECT 4.000 1063.200 1096.000 1065.880 ;
        RECT 4.400 1061.800 1096.000 1063.200 ;
        RECT 4.000 1057.760 1096.000 1061.800 ;
        RECT 4.000 1057.080 1095.600 1057.760 ;
        RECT 4.400 1056.360 1095.600 1057.080 ;
        RECT 4.400 1055.680 1096.000 1056.360 ;
        RECT 4.000 1050.960 1096.000 1055.680 ;
        RECT 4.400 1049.560 1096.000 1050.960 ;
        RECT 4.000 1048.240 1096.000 1049.560 ;
        RECT 4.000 1046.840 1095.600 1048.240 ;
        RECT 4.000 1045.520 1096.000 1046.840 ;
        RECT 4.400 1044.120 1096.000 1045.520 ;
        RECT 4.000 1039.400 1096.000 1044.120 ;
        RECT 4.400 1038.720 1096.000 1039.400 ;
        RECT 4.400 1038.000 1095.600 1038.720 ;
        RECT 4.000 1037.320 1095.600 1038.000 ;
        RECT 4.000 1033.960 1096.000 1037.320 ;
        RECT 4.400 1032.560 1096.000 1033.960 ;
        RECT 4.000 1029.200 1096.000 1032.560 ;
        RECT 4.000 1027.840 1095.600 1029.200 ;
        RECT 4.400 1027.800 1095.600 1027.840 ;
        RECT 4.400 1026.440 1096.000 1027.800 ;
        RECT 4.000 1022.400 1096.000 1026.440 ;
        RECT 4.400 1021.000 1096.000 1022.400 ;
        RECT 4.000 1019.680 1096.000 1021.000 ;
        RECT 4.000 1018.280 1095.600 1019.680 ;
        RECT 4.000 1016.280 1096.000 1018.280 ;
        RECT 4.400 1014.880 1096.000 1016.280 ;
        RECT 4.000 1010.840 1096.000 1014.880 ;
        RECT 4.400 1010.160 1096.000 1010.840 ;
        RECT 4.400 1009.440 1095.600 1010.160 ;
        RECT 4.000 1008.760 1095.600 1009.440 ;
        RECT 4.000 1004.720 1096.000 1008.760 ;
        RECT 4.400 1003.320 1096.000 1004.720 ;
        RECT 4.000 1000.640 1096.000 1003.320 ;
        RECT 4.000 999.240 1095.600 1000.640 ;
        RECT 4.000 998.600 1096.000 999.240 ;
        RECT 4.400 997.200 1096.000 998.600 ;
        RECT 4.000 993.160 1096.000 997.200 ;
        RECT 4.400 991.760 1096.000 993.160 ;
        RECT 4.000 991.120 1096.000 991.760 ;
        RECT 4.000 989.720 1095.600 991.120 ;
        RECT 4.000 987.040 1096.000 989.720 ;
        RECT 4.400 985.640 1096.000 987.040 ;
        RECT 4.000 981.600 1096.000 985.640 ;
        RECT 4.400 980.200 1095.600 981.600 ;
        RECT 4.000 975.480 1096.000 980.200 ;
        RECT 4.400 974.080 1096.000 975.480 ;
        RECT 4.000 972.080 1096.000 974.080 ;
        RECT 4.000 970.680 1095.600 972.080 ;
        RECT 4.000 970.040 1096.000 970.680 ;
        RECT 4.400 968.640 1096.000 970.040 ;
        RECT 4.000 963.920 1096.000 968.640 ;
        RECT 4.400 962.560 1096.000 963.920 ;
        RECT 4.400 962.520 1095.600 962.560 ;
        RECT 4.000 961.160 1095.600 962.520 ;
        RECT 4.000 957.800 1096.000 961.160 ;
        RECT 4.400 956.400 1096.000 957.800 ;
        RECT 4.000 953.040 1096.000 956.400 ;
        RECT 4.000 952.360 1095.600 953.040 ;
        RECT 4.400 951.640 1095.600 952.360 ;
        RECT 4.400 950.960 1096.000 951.640 ;
        RECT 4.000 946.240 1096.000 950.960 ;
        RECT 4.400 944.840 1096.000 946.240 ;
        RECT 4.000 943.520 1096.000 944.840 ;
        RECT 4.000 942.120 1095.600 943.520 ;
        RECT 4.000 940.800 1096.000 942.120 ;
        RECT 4.400 939.400 1096.000 940.800 ;
        RECT 4.000 934.680 1096.000 939.400 ;
        RECT 4.400 934.000 1096.000 934.680 ;
        RECT 4.400 933.280 1095.600 934.000 ;
        RECT 4.000 932.600 1095.600 933.280 ;
        RECT 4.000 929.240 1096.000 932.600 ;
        RECT 4.400 927.840 1096.000 929.240 ;
        RECT 4.000 924.480 1096.000 927.840 ;
        RECT 4.000 923.120 1095.600 924.480 ;
        RECT 4.400 923.080 1095.600 923.120 ;
        RECT 4.400 921.720 1096.000 923.080 ;
        RECT 4.000 917.680 1096.000 921.720 ;
        RECT 4.400 916.280 1096.000 917.680 ;
        RECT 4.000 915.640 1096.000 916.280 ;
        RECT 4.000 914.240 1095.600 915.640 ;
        RECT 4.000 911.560 1096.000 914.240 ;
        RECT 4.400 910.160 1096.000 911.560 ;
        RECT 4.000 906.120 1096.000 910.160 ;
        RECT 4.000 905.440 1095.600 906.120 ;
        RECT 4.400 904.720 1095.600 905.440 ;
        RECT 4.400 904.040 1096.000 904.720 ;
        RECT 4.000 900.000 1096.000 904.040 ;
        RECT 4.400 898.600 1096.000 900.000 ;
        RECT 4.000 896.600 1096.000 898.600 ;
        RECT 4.000 895.200 1095.600 896.600 ;
        RECT 4.000 893.880 1096.000 895.200 ;
        RECT 4.400 892.480 1096.000 893.880 ;
        RECT 4.000 888.440 1096.000 892.480 ;
        RECT 4.400 887.080 1096.000 888.440 ;
        RECT 4.400 887.040 1095.600 887.080 ;
        RECT 4.000 885.680 1095.600 887.040 ;
        RECT 4.000 882.320 1096.000 885.680 ;
        RECT 4.400 880.920 1096.000 882.320 ;
        RECT 4.000 877.560 1096.000 880.920 ;
        RECT 4.000 876.880 1095.600 877.560 ;
        RECT 4.400 876.160 1095.600 876.880 ;
        RECT 4.400 875.480 1096.000 876.160 ;
        RECT 4.000 870.760 1096.000 875.480 ;
        RECT 4.400 869.360 1096.000 870.760 ;
        RECT 4.000 868.040 1096.000 869.360 ;
        RECT 4.000 866.640 1095.600 868.040 ;
        RECT 4.000 865.320 1096.000 866.640 ;
        RECT 4.400 863.920 1096.000 865.320 ;
        RECT 4.000 859.200 1096.000 863.920 ;
        RECT 4.400 858.520 1096.000 859.200 ;
        RECT 4.400 857.800 1095.600 858.520 ;
        RECT 4.000 857.120 1095.600 857.800 ;
        RECT 4.000 853.080 1096.000 857.120 ;
        RECT 4.400 851.680 1096.000 853.080 ;
        RECT 4.000 849.000 1096.000 851.680 ;
        RECT 4.000 847.640 1095.600 849.000 ;
        RECT 4.400 847.600 1095.600 847.640 ;
        RECT 4.400 846.240 1096.000 847.600 ;
        RECT 4.000 841.520 1096.000 846.240 ;
        RECT 4.400 840.120 1096.000 841.520 ;
        RECT 4.000 839.480 1096.000 840.120 ;
        RECT 4.000 838.080 1095.600 839.480 ;
        RECT 4.000 836.080 1096.000 838.080 ;
        RECT 4.400 834.680 1096.000 836.080 ;
        RECT 4.000 829.960 1096.000 834.680 ;
        RECT 4.400 828.560 1095.600 829.960 ;
        RECT 4.000 824.520 1096.000 828.560 ;
        RECT 4.400 823.120 1096.000 824.520 ;
        RECT 4.000 820.440 1096.000 823.120 ;
        RECT 4.000 819.040 1095.600 820.440 ;
        RECT 4.000 818.400 1096.000 819.040 ;
        RECT 4.400 817.000 1096.000 818.400 ;
        RECT 4.000 812.280 1096.000 817.000 ;
        RECT 4.400 810.920 1096.000 812.280 ;
        RECT 4.400 810.880 1095.600 810.920 ;
        RECT 4.000 809.520 1095.600 810.880 ;
        RECT 4.000 806.840 1096.000 809.520 ;
        RECT 4.400 805.440 1096.000 806.840 ;
        RECT 4.000 801.400 1096.000 805.440 ;
        RECT 4.000 800.720 1095.600 801.400 ;
        RECT 4.400 800.000 1095.600 800.720 ;
        RECT 4.400 799.320 1096.000 800.000 ;
        RECT 4.000 795.280 1096.000 799.320 ;
        RECT 4.400 793.880 1096.000 795.280 ;
        RECT 4.000 791.880 1096.000 793.880 ;
        RECT 4.000 790.480 1095.600 791.880 ;
        RECT 4.000 789.160 1096.000 790.480 ;
        RECT 4.400 787.760 1096.000 789.160 ;
        RECT 4.000 783.720 1096.000 787.760 ;
        RECT 4.400 782.360 1096.000 783.720 ;
        RECT 4.400 782.320 1095.600 782.360 ;
        RECT 4.000 780.960 1095.600 782.320 ;
        RECT 4.000 777.600 1096.000 780.960 ;
        RECT 4.400 776.200 1096.000 777.600 ;
        RECT 4.000 772.840 1096.000 776.200 ;
        RECT 4.000 772.160 1095.600 772.840 ;
        RECT 4.400 771.440 1095.600 772.160 ;
        RECT 4.400 770.760 1096.000 771.440 ;
        RECT 4.000 766.040 1096.000 770.760 ;
        RECT 4.400 764.640 1096.000 766.040 ;
        RECT 4.000 763.320 1096.000 764.640 ;
        RECT 4.000 761.920 1095.600 763.320 ;
        RECT 4.000 759.920 1096.000 761.920 ;
        RECT 4.400 758.520 1096.000 759.920 ;
        RECT 4.000 754.480 1096.000 758.520 ;
        RECT 4.400 753.800 1096.000 754.480 ;
        RECT 4.400 753.080 1095.600 753.800 ;
        RECT 4.000 752.400 1095.600 753.080 ;
        RECT 4.000 748.360 1096.000 752.400 ;
        RECT 4.400 746.960 1096.000 748.360 ;
        RECT 4.000 744.280 1096.000 746.960 ;
        RECT 4.000 742.920 1095.600 744.280 ;
        RECT 4.400 742.880 1095.600 742.920 ;
        RECT 4.400 741.520 1096.000 742.880 ;
        RECT 4.000 736.800 1096.000 741.520 ;
        RECT 4.400 735.440 1096.000 736.800 ;
        RECT 4.400 735.400 1095.600 735.440 ;
        RECT 4.000 734.040 1095.600 735.400 ;
        RECT 4.000 731.360 1096.000 734.040 ;
        RECT 4.400 729.960 1096.000 731.360 ;
        RECT 4.000 725.920 1096.000 729.960 ;
        RECT 4.000 725.240 1095.600 725.920 ;
        RECT 4.400 724.520 1095.600 725.240 ;
        RECT 4.400 723.840 1096.000 724.520 ;
        RECT 4.000 719.120 1096.000 723.840 ;
        RECT 4.400 717.720 1096.000 719.120 ;
        RECT 4.000 716.400 1096.000 717.720 ;
        RECT 4.000 715.000 1095.600 716.400 ;
        RECT 4.000 713.680 1096.000 715.000 ;
        RECT 4.400 712.280 1096.000 713.680 ;
        RECT 4.000 707.560 1096.000 712.280 ;
        RECT 4.400 706.880 1096.000 707.560 ;
        RECT 4.400 706.160 1095.600 706.880 ;
        RECT 4.000 705.480 1095.600 706.160 ;
        RECT 4.000 702.120 1096.000 705.480 ;
        RECT 4.400 700.720 1096.000 702.120 ;
        RECT 4.000 697.360 1096.000 700.720 ;
        RECT 4.000 696.000 1095.600 697.360 ;
        RECT 4.400 695.960 1095.600 696.000 ;
        RECT 4.400 694.600 1096.000 695.960 ;
        RECT 4.000 690.560 1096.000 694.600 ;
        RECT 4.400 689.160 1096.000 690.560 ;
        RECT 4.000 687.840 1096.000 689.160 ;
        RECT 4.000 686.440 1095.600 687.840 ;
        RECT 4.000 684.440 1096.000 686.440 ;
        RECT 4.400 683.040 1096.000 684.440 ;
        RECT 4.000 679.000 1096.000 683.040 ;
        RECT 4.400 678.320 1096.000 679.000 ;
        RECT 4.400 677.600 1095.600 678.320 ;
        RECT 4.000 676.920 1095.600 677.600 ;
        RECT 4.000 672.880 1096.000 676.920 ;
        RECT 4.400 671.480 1096.000 672.880 ;
        RECT 4.000 668.800 1096.000 671.480 ;
        RECT 4.000 667.400 1095.600 668.800 ;
        RECT 4.000 666.760 1096.000 667.400 ;
        RECT 4.400 665.360 1096.000 666.760 ;
        RECT 4.000 661.320 1096.000 665.360 ;
        RECT 4.400 659.920 1096.000 661.320 ;
        RECT 4.000 659.280 1096.000 659.920 ;
        RECT 4.000 657.880 1095.600 659.280 ;
        RECT 4.000 655.200 1096.000 657.880 ;
        RECT 4.400 653.800 1096.000 655.200 ;
        RECT 4.000 649.760 1096.000 653.800 ;
        RECT 4.400 648.360 1095.600 649.760 ;
        RECT 4.000 643.640 1096.000 648.360 ;
        RECT 4.400 642.240 1096.000 643.640 ;
        RECT 4.000 640.240 1096.000 642.240 ;
        RECT 4.000 638.840 1095.600 640.240 ;
        RECT 4.000 638.200 1096.000 638.840 ;
        RECT 4.400 636.800 1096.000 638.200 ;
        RECT 4.000 632.080 1096.000 636.800 ;
        RECT 4.400 630.720 1096.000 632.080 ;
        RECT 4.400 630.680 1095.600 630.720 ;
        RECT 4.000 629.320 1095.600 630.680 ;
        RECT 4.000 626.640 1096.000 629.320 ;
        RECT 4.400 625.240 1096.000 626.640 ;
        RECT 4.000 621.200 1096.000 625.240 ;
        RECT 4.000 620.520 1095.600 621.200 ;
        RECT 4.400 619.800 1095.600 620.520 ;
        RECT 4.400 619.120 1096.000 619.800 ;
        RECT 4.000 614.400 1096.000 619.120 ;
        RECT 4.400 613.000 1096.000 614.400 ;
        RECT 4.000 611.680 1096.000 613.000 ;
        RECT 4.000 610.280 1095.600 611.680 ;
        RECT 4.000 608.960 1096.000 610.280 ;
        RECT 4.400 607.560 1096.000 608.960 ;
        RECT 4.000 602.840 1096.000 607.560 ;
        RECT 4.400 602.160 1096.000 602.840 ;
        RECT 4.400 601.440 1095.600 602.160 ;
        RECT 4.000 600.760 1095.600 601.440 ;
        RECT 4.000 597.400 1096.000 600.760 ;
        RECT 4.400 596.000 1096.000 597.400 ;
        RECT 4.000 592.640 1096.000 596.000 ;
        RECT 4.000 591.280 1095.600 592.640 ;
        RECT 4.400 591.240 1095.600 591.280 ;
        RECT 4.400 589.880 1096.000 591.240 ;
        RECT 4.000 585.840 1096.000 589.880 ;
        RECT 4.400 584.440 1096.000 585.840 ;
        RECT 4.000 583.120 1096.000 584.440 ;
        RECT 4.000 581.720 1095.600 583.120 ;
        RECT 4.000 579.720 1096.000 581.720 ;
        RECT 4.400 578.320 1096.000 579.720 ;
        RECT 4.000 573.600 1096.000 578.320 ;
        RECT 4.400 572.200 1095.600 573.600 ;
        RECT 4.000 568.160 1096.000 572.200 ;
        RECT 4.400 566.760 1096.000 568.160 ;
        RECT 4.000 564.080 1096.000 566.760 ;
        RECT 4.000 562.680 1095.600 564.080 ;
        RECT 4.000 562.040 1096.000 562.680 ;
        RECT 4.400 560.640 1096.000 562.040 ;
        RECT 4.000 556.600 1096.000 560.640 ;
        RECT 4.400 555.240 1096.000 556.600 ;
        RECT 4.400 555.200 1095.600 555.240 ;
        RECT 4.000 553.840 1095.600 555.200 ;
        RECT 4.000 550.480 1096.000 553.840 ;
        RECT 4.400 549.080 1096.000 550.480 ;
        RECT 4.000 545.720 1096.000 549.080 ;
        RECT 4.000 545.040 1095.600 545.720 ;
        RECT 4.400 544.320 1095.600 545.040 ;
        RECT 4.400 543.640 1096.000 544.320 ;
        RECT 4.000 538.920 1096.000 543.640 ;
        RECT 4.400 537.520 1096.000 538.920 ;
        RECT 4.000 536.200 1096.000 537.520 ;
        RECT 4.000 534.800 1095.600 536.200 ;
        RECT 4.000 533.480 1096.000 534.800 ;
        RECT 4.400 532.080 1096.000 533.480 ;
        RECT 4.000 527.360 1096.000 532.080 ;
        RECT 4.400 526.680 1096.000 527.360 ;
        RECT 4.400 525.960 1095.600 526.680 ;
        RECT 4.000 525.280 1095.600 525.960 ;
        RECT 4.000 521.240 1096.000 525.280 ;
        RECT 4.400 519.840 1096.000 521.240 ;
        RECT 4.000 517.160 1096.000 519.840 ;
        RECT 4.000 515.800 1095.600 517.160 ;
        RECT 4.400 515.760 1095.600 515.800 ;
        RECT 4.400 514.400 1096.000 515.760 ;
        RECT 4.000 509.680 1096.000 514.400 ;
        RECT 4.400 508.280 1096.000 509.680 ;
        RECT 4.000 507.640 1096.000 508.280 ;
        RECT 4.000 506.240 1095.600 507.640 ;
        RECT 4.000 504.240 1096.000 506.240 ;
        RECT 4.400 502.840 1096.000 504.240 ;
        RECT 4.000 498.120 1096.000 502.840 ;
        RECT 4.400 496.720 1095.600 498.120 ;
        RECT 4.000 492.680 1096.000 496.720 ;
        RECT 4.400 491.280 1096.000 492.680 ;
        RECT 4.000 488.600 1096.000 491.280 ;
        RECT 4.000 487.200 1095.600 488.600 ;
        RECT 4.000 486.560 1096.000 487.200 ;
        RECT 4.400 485.160 1096.000 486.560 ;
        RECT 4.000 480.440 1096.000 485.160 ;
        RECT 4.400 479.080 1096.000 480.440 ;
        RECT 4.400 479.040 1095.600 479.080 ;
        RECT 4.000 477.680 1095.600 479.040 ;
        RECT 4.000 475.000 1096.000 477.680 ;
        RECT 4.400 473.600 1096.000 475.000 ;
        RECT 4.000 469.560 1096.000 473.600 ;
        RECT 4.000 468.880 1095.600 469.560 ;
        RECT 4.400 468.160 1095.600 468.880 ;
        RECT 4.400 467.480 1096.000 468.160 ;
        RECT 4.000 463.440 1096.000 467.480 ;
        RECT 4.400 462.040 1096.000 463.440 ;
        RECT 4.000 460.040 1096.000 462.040 ;
        RECT 4.000 458.640 1095.600 460.040 ;
        RECT 4.000 457.320 1096.000 458.640 ;
        RECT 4.400 455.920 1096.000 457.320 ;
        RECT 4.000 451.880 1096.000 455.920 ;
        RECT 4.400 450.520 1096.000 451.880 ;
        RECT 4.400 450.480 1095.600 450.520 ;
        RECT 4.000 449.120 1095.600 450.480 ;
        RECT 4.000 445.760 1096.000 449.120 ;
        RECT 4.400 444.360 1096.000 445.760 ;
        RECT 4.000 441.000 1096.000 444.360 ;
        RECT 4.000 440.320 1095.600 441.000 ;
        RECT 4.400 439.600 1095.600 440.320 ;
        RECT 4.400 438.920 1096.000 439.600 ;
        RECT 4.000 434.200 1096.000 438.920 ;
        RECT 4.400 432.800 1096.000 434.200 ;
        RECT 4.000 431.480 1096.000 432.800 ;
        RECT 4.000 430.080 1095.600 431.480 ;
        RECT 4.000 428.080 1096.000 430.080 ;
        RECT 4.400 426.680 1096.000 428.080 ;
        RECT 4.000 422.640 1096.000 426.680 ;
        RECT 4.400 421.960 1096.000 422.640 ;
        RECT 4.400 421.240 1095.600 421.960 ;
        RECT 4.000 420.560 1095.600 421.240 ;
        RECT 4.000 416.520 1096.000 420.560 ;
        RECT 4.400 415.120 1096.000 416.520 ;
        RECT 4.000 412.440 1096.000 415.120 ;
        RECT 4.000 411.080 1095.600 412.440 ;
        RECT 4.400 411.040 1095.600 411.080 ;
        RECT 4.400 409.680 1096.000 411.040 ;
        RECT 4.000 404.960 1096.000 409.680 ;
        RECT 4.400 403.560 1096.000 404.960 ;
        RECT 4.000 402.920 1096.000 403.560 ;
        RECT 4.000 401.520 1095.600 402.920 ;
        RECT 4.000 399.520 1096.000 401.520 ;
        RECT 4.400 398.120 1096.000 399.520 ;
        RECT 4.000 393.400 1096.000 398.120 ;
        RECT 4.400 392.000 1095.600 393.400 ;
        RECT 4.000 387.960 1096.000 392.000 ;
        RECT 4.400 386.560 1096.000 387.960 ;
        RECT 4.000 383.880 1096.000 386.560 ;
        RECT 4.000 382.480 1095.600 383.880 ;
        RECT 4.000 381.840 1096.000 382.480 ;
        RECT 4.400 380.440 1096.000 381.840 ;
        RECT 4.000 375.720 1096.000 380.440 ;
        RECT 4.400 374.360 1096.000 375.720 ;
        RECT 4.400 374.320 1095.600 374.360 ;
        RECT 4.000 372.960 1095.600 374.320 ;
        RECT 4.000 370.280 1096.000 372.960 ;
        RECT 4.400 368.880 1096.000 370.280 ;
        RECT 4.000 365.520 1096.000 368.880 ;
        RECT 4.000 364.160 1095.600 365.520 ;
        RECT 4.400 364.120 1095.600 364.160 ;
        RECT 4.400 362.760 1096.000 364.120 ;
        RECT 4.000 358.720 1096.000 362.760 ;
        RECT 4.400 357.320 1096.000 358.720 ;
        RECT 4.000 356.000 1096.000 357.320 ;
        RECT 4.000 354.600 1095.600 356.000 ;
        RECT 4.000 352.600 1096.000 354.600 ;
        RECT 4.400 351.200 1096.000 352.600 ;
        RECT 4.000 347.160 1096.000 351.200 ;
        RECT 4.400 346.480 1096.000 347.160 ;
        RECT 4.400 345.760 1095.600 346.480 ;
        RECT 4.000 345.080 1095.600 345.760 ;
        RECT 4.000 341.040 1096.000 345.080 ;
        RECT 4.400 339.640 1096.000 341.040 ;
        RECT 4.000 336.960 1096.000 339.640 ;
        RECT 4.000 335.560 1095.600 336.960 ;
        RECT 4.000 334.920 1096.000 335.560 ;
        RECT 4.400 333.520 1096.000 334.920 ;
        RECT 4.000 329.480 1096.000 333.520 ;
        RECT 4.400 328.080 1096.000 329.480 ;
        RECT 4.000 327.440 1096.000 328.080 ;
        RECT 4.000 326.040 1095.600 327.440 ;
        RECT 4.000 323.360 1096.000 326.040 ;
        RECT 4.400 321.960 1096.000 323.360 ;
        RECT 4.000 317.920 1096.000 321.960 ;
        RECT 4.400 316.520 1095.600 317.920 ;
        RECT 4.000 311.800 1096.000 316.520 ;
        RECT 4.400 310.400 1096.000 311.800 ;
        RECT 4.000 308.400 1096.000 310.400 ;
        RECT 4.000 307.000 1095.600 308.400 ;
        RECT 4.000 306.360 1096.000 307.000 ;
        RECT 4.400 304.960 1096.000 306.360 ;
        RECT 4.000 300.240 1096.000 304.960 ;
        RECT 4.400 298.880 1096.000 300.240 ;
        RECT 4.400 298.840 1095.600 298.880 ;
        RECT 4.000 297.480 1095.600 298.840 ;
        RECT 4.000 294.800 1096.000 297.480 ;
        RECT 4.400 293.400 1096.000 294.800 ;
        RECT 4.000 289.360 1096.000 293.400 ;
        RECT 4.000 288.680 1095.600 289.360 ;
        RECT 4.400 287.960 1095.600 288.680 ;
        RECT 4.400 287.280 1096.000 287.960 ;
        RECT 4.000 282.560 1096.000 287.280 ;
        RECT 4.400 281.160 1096.000 282.560 ;
        RECT 4.000 279.840 1096.000 281.160 ;
        RECT 4.000 278.440 1095.600 279.840 ;
        RECT 4.000 277.120 1096.000 278.440 ;
        RECT 4.400 275.720 1096.000 277.120 ;
        RECT 4.000 271.000 1096.000 275.720 ;
        RECT 4.400 270.320 1096.000 271.000 ;
        RECT 4.400 269.600 1095.600 270.320 ;
        RECT 4.000 268.920 1095.600 269.600 ;
        RECT 4.000 265.560 1096.000 268.920 ;
        RECT 4.400 264.160 1096.000 265.560 ;
        RECT 4.000 260.800 1096.000 264.160 ;
        RECT 4.000 259.440 1095.600 260.800 ;
        RECT 4.400 259.400 1095.600 259.440 ;
        RECT 4.400 258.040 1096.000 259.400 ;
        RECT 4.000 254.000 1096.000 258.040 ;
        RECT 4.400 252.600 1096.000 254.000 ;
        RECT 4.000 251.280 1096.000 252.600 ;
        RECT 4.000 249.880 1095.600 251.280 ;
        RECT 4.000 247.880 1096.000 249.880 ;
        RECT 4.400 246.480 1096.000 247.880 ;
        RECT 4.000 241.760 1096.000 246.480 ;
        RECT 4.400 240.360 1095.600 241.760 ;
        RECT 4.000 236.320 1096.000 240.360 ;
        RECT 4.400 234.920 1096.000 236.320 ;
        RECT 4.000 232.240 1096.000 234.920 ;
        RECT 4.000 230.840 1095.600 232.240 ;
        RECT 4.000 230.200 1096.000 230.840 ;
        RECT 4.400 228.800 1096.000 230.200 ;
        RECT 4.000 224.760 1096.000 228.800 ;
        RECT 4.400 223.360 1096.000 224.760 ;
        RECT 4.000 222.720 1096.000 223.360 ;
        RECT 4.000 221.320 1095.600 222.720 ;
        RECT 4.000 218.640 1096.000 221.320 ;
        RECT 4.400 217.240 1096.000 218.640 ;
        RECT 4.000 213.200 1096.000 217.240 ;
        RECT 4.400 211.800 1095.600 213.200 ;
        RECT 4.000 207.080 1096.000 211.800 ;
        RECT 4.400 205.680 1096.000 207.080 ;
        RECT 4.000 203.680 1096.000 205.680 ;
        RECT 4.000 202.280 1095.600 203.680 ;
        RECT 4.000 201.640 1096.000 202.280 ;
        RECT 4.400 200.240 1096.000 201.640 ;
        RECT 4.000 195.520 1096.000 200.240 ;
        RECT 4.400 194.160 1096.000 195.520 ;
        RECT 4.400 194.120 1095.600 194.160 ;
        RECT 4.000 192.760 1095.600 194.120 ;
        RECT 4.000 189.400 1096.000 192.760 ;
        RECT 4.400 188.000 1096.000 189.400 ;
        RECT 4.000 185.320 1096.000 188.000 ;
        RECT 4.000 183.960 1095.600 185.320 ;
        RECT 4.400 183.920 1095.600 183.960 ;
        RECT 4.400 182.560 1096.000 183.920 ;
        RECT 4.000 177.840 1096.000 182.560 ;
        RECT 4.400 176.440 1096.000 177.840 ;
        RECT 4.000 175.800 1096.000 176.440 ;
        RECT 4.000 174.400 1095.600 175.800 ;
        RECT 4.000 172.400 1096.000 174.400 ;
        RECT 4.400 171.000 1096.000 172.400 ;
        RECT 4.000 166.280 1096.000 171.000 ;
        RECT 4.400 164.880 1095.600 166.280 ;
        RECT 4.000 160.840 1096.000 164.880 ;
        RECT 4.400 159.440 1096.000 160.840 ;
        RECT 4.000 156.760 1096.000 159.440 ;
        RECT 4.000 155.360 1095.600 156.760 ;
        RECT 4.000 154.720 1096.000 155.360 ;
        RECT 4.400 153.320 1096.000 154.720 ;
        RECT 4.000 149.280 1096.000 153.320 ;
        RECT 4.400 147.880 1096.000 149.280 ;
        RECT 4.000 147.240 1096.000 147.880 ;
        RECT 4.000 145.840 1095.600 147.240 ;
        RECT 4.000 143.160 1096.000 145.840 ;
        RECT 4.400 141.760 1096.000 143.160 ;
        RECT 4.000 137.720 1096.000 141.760 ;
        RECT 4.000 137.040 1095.600 137.720 ;
        RECT 4.400 136.320 1095.600 137.040 ;
        RECT 4.400 135.640 1096.000 136.320 ;
        RECT 4.000 131.600 1096.000 135.640 ;
        RECT 4.400 130.200 1096.000 131.600 ;
        RECT 4.000 128.200 1096.000 130.200 ;
        RECT 4.000 126.800 1095.600 128.200 ;
        RECT 4.000 125.480 1096.000 126.800 ;
        RECT 4.400 124.080 1096.000 125.480 ;
        RECT 4.000 120.040 1096.000 124.080 ;
        RECT 4.400 118.680 1096.000 120.040 ;
        RECT 4.400 118.640 1095.600 118.680 ;
        RECT 4.000 117.280 1095.600 118.640 ;
        RECT 4.000 113.920 1096.000 117.280 ;
        RECT 4.400 112.520 1096.000 113.920 ;
        RECT 4.000 109.160 1096.000 112.520 ;
        RECT 4.000 108.480 1095.600 109.160 ;
        RECT 4.400 107.760 1095.600 108.480 ;
        RECT 4.400 107.080 1096.000 107.760 ;
        RECT 4.000 102.360 1096.000 107.080 ;
        RECT 4.400 100.960 1096.000 102.360 ;
        RECT 4.000 99.640 1096.000 100.960 ;
        RECT 4.000 98.240 1095.600 99.640 ;
        RECT 4.000 96.240 1096.000 98.240 ;
        RECT 4.400 94.840 1096.000 96.240 ;
        RECT 4.000 90.800 1096.000 94.840 ;
        RECT 4.400 90.120 1096.000 90.800 ;
        RECT 4.400 89.400 1095.600 90.120 ;
        RECT 4.000 88.720 1095.600 89.400 ;
        RECT 4.000 84.680 1096.000 88.720 ;
        RECT 4.400 83.280 1096.000 84.680 ;
        RECT 4.000 80.600 1096.000 83.280 ;
        RECT 4.000 79.240 1095.600 80.600 ;
        RECT 4.400 79.200 1095.600 79.240 ;
        RECT 4.400 77.840 1096.000 79.200 ;
        RECT 4.000 73.120 1096.000 77.840 ;
        RECT 4.400 71.720 1096.000 73.120 ;
        RECT 4.000 71.080 1096.000 71.720 ;
        RECT 4.000 69.680 1095.600 71.080 ;
        RECT 4.000 67.680 1096.000 69.680 ;
        RECT 4.400 66.280 1096.000 67.680 ;
        RECT 4.000 61.560 1096.000 66.280 ;
        RECT 4.400 60.160 1095.600 61.560 ;
        RECT 4.000 56.120 1096.000 60.160 ;
        RECT 4.400 54.720 1096.000 56.120 ;
        RECT 4.000 52.040 1096.000 54.720 ;
        RECT 4.000 50.640 1095.600 52.040 ;
        RECT 4.000 50.000 1096.000 50.640 ;
        RECT 4.400 48.600 1096.000 50.000 ;
        RECT 4.000 43.880 1096.000 48.600 ;
        RECT 4.400 42.520 1096.000 43.880 ;
        RECT 4.400 42.480 1095.600 42.520 ;
        RECT 4.000 41.120 1095.600 42.480 ;
        RECT 4.000 38.440 1096.000 41.120 ;
        RECT 4.400 37.040 1096.000 38.440 ;
        RECT 4.000 33.000 1096.000 37.040 ;
        RECT 4.000 32.320 1095.600 33.000 ;
        RECT 4.400 31.600 1095.600 32.320 ;
        RECT 4.400 30.920 1096.000 31.600 ;
        RECT 4.000 26.880 1096.000 30.920 ;
        RECT 4.400 25.480 1096.000 26.880 ;
        RECT 4.000 23.480 1096.000 25.480 ;
        RECT 4.000 22.080 1095.600 23.480 ;
        RECT 4.000 20.760 1096.000 22.080 ;
        RECT 4.400 19.360 1096.000 20.760 ;
        RECT 4.000 15.320 1096.000 19.360 ;
        RECT 4.400 13.960 1096.000 15.320 ;
        RECT 4.400 13.920 1095.600 13.960 ;
        RECT 4.000 12.560 1095.600 13.920 ;
        RECT 4.000 9.200 1096.000 12.560 ;
        RECT 4.400 7.800 1096.000 9.200 ;
        RECT 4.000 5.120 1096.000 7.800 ;
        RECT 4.000 3.760 1095.600 5.120 ;
        RECT 4.400 3.720 1095.600 3.760 ;
        RECT 4.400 2.895 1096.000 3.720 ;
      LAYER met4 ;
        RECT 10.415 12.415 20.640 1086.465 ;
        RECT 23.040 12.415 97.440 1086.465 ;
        RECT 99.840 12.415 174.240 1086.465 ;
        RECT 176.640 12.415 251.040 1086.465 ;
        RECT 253.440 12.415 327.840 1086.465 ;
        RECT 330.240 12.415 404.640 1086.465 ;
        RECT 407.040 12.415 481.440 1086.465 ;
        RECT 483.840 12.415 558.240 1086.465 ;
        RECT 560.640 12.415 635.040 1086.465 ;
        RECT 637.440 12.415 711.840 1086.465 ;
        RECT 714.240 12.415 788.640 1086.465 ;
        RECT 791.040 12.415 865.440 1086.465 ;
        RECT 867.840 12.415 942.240 1086.465 ;
        RECT 944.640 12.415 1019.040 1086.465 ;
        RECT 1021.440 12.415 1088.985 1086.465 ;
  END
END WB_InterConnect
END LIBRARY

