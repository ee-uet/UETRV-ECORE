magic
tech sky130A
magscale 1 2
timestamp 1647757248
<< obsli1 >>
rect 1104 2159 98808 97393
<< obsm1 >>
rect 1104 2128 98808 97424
<< metal2 >>
rect 2778 99200 2834 100000
rect 8298 99200 8354 100000
rect 13818 99200 13874 100000
rect 19430 99200 19486 100000
rect 24950 99200 25006 100000
rect 30470 99200 30526 100000
rect 36082 99200 36138 100000
rect 41602 99200 41658 100000
rect 47214 99200 47270 100000
rect 52734 99200 52790 100000
rect 58254 99200 58310 100000
rect 63866 99200 63922 100000
rect 69386 99200 69442 100000
rect 74998 99200 75054 100000
rect 80518 99200 80574 100000
rect 86038 99200 86094 100000
rect 91650 99200 91706 100000
rect 97170 99200 97226 100000
rect 1766 0 1822 800
rect 5262 0 5318 800
rect 8850 0 8906 800
rect 12438 0 12494 800
rect 16026 0 16082 800
rect 19614 0 19670 800
rect 23110 0 23166 800
rect 26698 0 26754 800
rect 30286 0 30342 800
rect 33874 0 33930 800
rect 37462 0 37518 800
rect 41050 0 41106 800
rect 44546 0 44602 800
rect 48134 0 48190 800
rect 51722 0 51778 800
rect 55310 0 55366 800
rect 58898 0 58954 800
rect 62394 0 62450 800
rect 65982 0 66038 800
rect 69570 0 69626 800
rect 73158 0 73214 800
rect 76746 0 76802 800
rect 80334 0 80390 800
rect 83830 0 83886 800
rect 87418 0 87474 800
rect 91006 0 91062 800
rect 94594 0 94650 800
rect 98182 0 98238 800
<< obsm2 >>
rect 1398 99144 2722 99362
rect 2890 99144 8242 99362
rect 8410 99144 13762 99362
rect 13930 99144 19374 99362
rect 19542 99144 24894 99362
rect 25062 99144 30414 99362
rect 30582 99144 36026 99362
rect 36194 99144 41546 99362
rect 41714 99144 47158 99362
rect 47326 99144 52678 99362
rect 52846 99144 58198 99362
rect 58366 99144 63810 99362
rect 63978 99144 69330 99362
rect 69498 99144 74942 99362
rect 75110 99144 80462 99362
rect 80630 99144 85982 99362
rect 86150 99144 91594 99362
rect 91762 99144 97114 99362
rect 97282 99144 98330 99362
rect 1398 856 98330 99144
rect 1398 734 1710 856
rect 1878 734 5206 856
rect 5374 734 8794 856
rect 8962 734 12382 856
rect 12550 734 15970 856
rect 16138 734 19558 856
rect 19726 734 23054 856
rect 23222 734 26642 856
rect 26810 734 30230 856
rect 30398 734 33818 856
rect 33986 734 37406 856
rect 37574 734 40994 856
rect 41162 734 44490 856
rect 44658 734 48078 856
rect 48246 734 51666 856
rect 51834 734 55254 856
rect 55422 734 58842 856
rect 59010 734 62338 856
rect 62506 734 65926 856
rect 66094 734 69514 856
rect 69682 734 73102 856
rect 73270 734 76690 856
rect 76858 734 80278 856
rect 80446 734 83774 856
rect 83942 734 87362 856
rect 87530 734 90950 856
rect 91118 734 94538 856
rect 94706 734 98126 856
rect 98294 734 98330 856
<< metal3 >>
rect 0 97928 800 98048
rect 99200 97520 100000 97640
rect 0 94256 800 94376
rect 99200 93032 100000 93152
rect 0 90584 800 90704
rect 99200 88408 100000 88528
rect 0 86912 800 87032
rect 99200 83920 100000 84040
rect 0 83104 800 83224
rect 0 79432 800 79552
rect 99200 79296 100000 79416
rect 0 75760 800 75880
rect 99200 74808 100000 74928
rect 0 72088 800 72208
rect 99200 70320 100000 70440
rect 0 68416 800 68536
rect 99200 65696 100000 65816
rect 0 64608 800 64728
rect 99200 61208 100000 61328
rect 0 60936 800 61056
rect 0 57264 800 57384
rect 99200 56584 100000 56704
rect 0 53592 800 53712
rect 99200 52096 100000 52216
rect 0 49784 800 49904
rect 99200 47608 100000 47728
rect 0 46112 800 46232
rect 99200 42984 100000 43104
rect 0 42440 800 42560
rect 0 38768 800 38888
rect 99200 38496 100000 38616
rect 0 35096 800 35216
rect 99200 33872 100000 33992
rect 0 31288 800 31408
rect 99200 29384 100000 29504
rect 0 27616 800 27736
rect 99200 24896 100000 25016
rect 0 23944 800 24064
rect 0 20272 800 20392
rect 99200 20272 100000 20392
rect 0 16464 800 16584
rect 99200 15784 100000 15904
rect 0 12792 800 12912
rect 99200 11160 100000 11280
rect 0 9120 800 9240
rect 99200 6672 100000 6792
rect 0 5448 800 5568
rect 99200 2184 100000 2304
rect 0 1776 800 1896
<< obsm3 >>
rect 880 97848 99200 98021
rect 800 97720 99200 97848
rect 800 97440 99120 97720
rect 800 94456 99200 97440
rect 880 94176 99200 94456
rect 800 93232 99200 94176
rect 800 92952 99120 93232
rect 800 90784 99200 92952
rect 880 90504 99200 90784
rect 800 88608 99200 90504
rect 800 88328 99120 88608
rect 800 87112 99200 88328
rect 880 86832 99200 87112
rect 800 84120 99200 86832
rect 800 83840 99120 84120
rect 800 83304 99200 83840
rect 880 83024 99200 83304
rect 800 79632 99200 83024
rect 880 79496 99200 79632
rect 880 79352 99120 79496
rect 800 79216 99120 79352
rect 800 75960 99200 79216
rect 880 75680 99200 75960
rect 800 75008 99200 75680
rect 800 74728 99120 75008
rect 800 72288 99200 74728
rect 880 72008 99200 72288
rect 800 70520 99200 72008
rect 800 70240 99120 70520
rect 800 68616 99200 70240
rect 880 68336 99200 68616
rect 800 65896 99200 68336
rect 800 65616 99120 65896
rect 800 64808 99200 65616
rect 880 64528 99200 64808
rect 800 61408 99200 64528
rect 800 61136 99120 61408
rect 880 61128 99120 61136
rect 880 60856 99200 61128
rect 800 57464 99200 60856
rect 880 57184 99200 57464
rect 800 56784 99200 57184
rect 800 56504 99120 56784
rect 800 53792 99200 56504
rect 880 53512 99200 53792
rect 800 52296 99200 53512
rect 800 52016 99120 52296
rect 800 49984 99200 52016
rect 880 49704 99200 49984
rect 800 47808 99200 49704
rect 800 47528 99120 47808
rect 800 46312 99200 47528
rect 880 46032 99200 46312
rect 800 43184 99200 46032
rect 800 42904 99120 43184
rect 800 42640 99200 42904
rect 880 42360 99200 42640
rect 800 38968 99200 42360
rect 880 38696 99200 38968
rect 880 38688 99120 38696
rect 800 38416 99120 38688
rect 800 35296 99200 38416
rect 880 35016 99200 35296
rect 800 34072 99200 35016
rect 800 33792 99120 34072
rect 800 31488 99200 33792
rect 880 31208 99200 31488
rect 800 29584 99200 31208
rect 800 29304 99120 29584
rect 800 27816 99200 29304
rect 880 27536 99200 27816
rect 800 25096 99200 27536
rect 800 24816 99120 25096
rect 800 24144 99200 24816
rect 880 23864 99200 24144
rect 800 20472 99200 23864
rect 880 20192 99120 20472
rect 800 16664 99200 20192
rect 880 16384 99200 16664
rect 800 15984 99200 16384
rect 800 15704 99120 15984
rect 800 12992 99200 15704
rect 880 12712 99200 12992
rect 800 11360 99200 12712
rect 800 11080 99120 11360
rect 800 9320 99200 11080
rect 880 9040 99200 9320
rect 800 6872 99200 9040
rect 800 6592 99120 6872
rect 800 5648 99200 6592
rect 880 5368 99200 5648
rect 800 2384 99200 5368
rect 800 2104 99120 2384
rect 800 1976 99200 2104
rect 880 1803 99200 1976
<< metal4 >>
rect 4208 2128 4528 97424
rect 19568 2128 19888 97424
rect 34928 2128 35248 97424
rect 50288 2128 50608 97424
rect 65648 2128 65968 97424
rect 81008 2128 81328 97424
rect 96368 2128 96688 97424
<< obsm4 >>
rect 13491 2211 19488 96661
rect 19968 2211 34848 96661
rect 35328 2211 50208 96661
rect 50688 2211 65568 96661
rect 66048 2211 80928 96661
rect 81408 2211 87157 96661
<< labels >>
rlabel metal2 s 1766 0 1822 800 6 clock
port 1 nsew signal input
rlabel metal3 s 99200 2184 100000 2304 6 io_ba_match
port 2 nsew signal input
rlabel metal3 s 0 1776 800 1896 6 io_motor_irq
port 3 nsew signal output
rlabel metal2 s 2778 99200 2834 100000 6 io_pwm_high
port 4 nsew signal output
rlabel metal2 s 8298 99200 8354 100000 6 io_pwm_low
port 5 nsew signal output
rlabel metal3 s 99200 6672 100000 6792 6 io_qei_ch_a
port 6 nsew signal input
rlabel metal2 s 8850 0 8906 800 6 io_qei_ch_b
port 7 nsew signal input
rlabel metal3 s 0 5448 800 5568 6 io_wbs_ack_o
port 8 nsew signal output
rlabel metal2 s 13818 99200 13874 100000 6 io_wbs_data_o[0]
port 9 nsew signal output
rlabel metal2 s 58254 99200 58310 100000 6 io_wbs_data_o[10]
port 10 nsew signal output
rlabel metal2 s 55310 0 55366 800 6 io_wbs_data_o[11]
port 11 nsew signal output
rlabel metal3 s 0 38768 800 38888 6 io_wbs_data_o[12]
port 12 nsew signal output
rlabel metal2 s 65982 0 66038 800 6 io_wbs_data_o[13]
port 13 nsew signal output
rlabel metal3 s 99200 65696 100000 65816 6 io_wbs_data_o[14]
port 14 nsew signal output
rlabel metal3 s 99200 74808 100000 74928 6 io_wbs_data_o[15]
port 15 nsew signal output
rlabel metal2 s 76746 0 76802 800 6 io_wbs_data_o[16]
port 16 nsew signal output
rlabel metal3 s 0 46112 800 46232 6 io_wbs_data_o[17]
port 17 nsew signal output
rlabel metal2 s 83830 0 83886 800 6 io_wbs_data_o[18]
port 18 nsew signal output
rlabel metal3 s 0 53592 800 53712 6 io_wbs_data_o[19]
port 19 nsew signal output
rlabel metal3 s 0 12792 800 12912 6 io_wbs_data_o[1]
port 20 nsew signal output
rlabel metal3 s 99200 79296 100000 79416 6 io_wbs_data_o[20]
port 21 nsew signal output
rlabel metal3 s 0 60936 800 61056 6 io_wbs_data_o[21]
port 22 nsew signal output
rlabel metal2 s 80518 99200 80574 100000 6 io_wbs_data_o[22]
port 23 nsew signal output
rlabel metal3 s 99200 83920 100000 84040 6 io_wbs_data_o[23]
port 24 nsew signal output
rlabel metal3 s 99200 93032 100000 93152 6 io_wbs_data_o[24]
port 25 nsew signal output
rlabel metal2 s 91006 0 91062 800 6 io_wbs_data_o[25]
port 26 nsew signal output
rlabel metal3 s 0 72088 800 72208 6 io_wbs_data_o[26]
port 27 nsew signal output
rlabel metal3 s 0 79432 800 79552 6 io_wbs_data_o[27]
port 28 nsew signal output
rlabel metal3 s 0 86912 800 87032 6 io_wbs_data_o[28]
port 29 nsew signal output
rlabel metal2 s 94594 0 94650 800 6 io_wbs_data_o[29]
port 30 nsew signal output
rlabel metal3 s 99200 29384 100000 29504 6 io_wbs_data_o[2]
port 31 nsew signal output
rlabel metal3 s 0 94256 800 94376 6 io_wbs_data_o[30]
port 32 nsew signal output
rlabel metal2 s 97170 99200 97226 100000 6 io_wbs_data_o[31]
port 33 nsew signal output
rlabel metal2 s 19614 0 19670 800 6 io_wbs_data_o[3]
port 34 nsew signal output
rlabel metal2 s 23110 0 23166 800 6 io_wbs_data_o[4]
port 35 nsew signal output
rlabel metal3 s 99200 42984 100000 43104 6 io_wbs_data_o[5]
port 36 nsew signal output
rlabel metal3 s 99200 47608 100000 47728 6 io_wbs_data_o[6]
port 37 nsew signal output
rlabel metal3 s 0 27616 800 27736 6 io_wbs_data_o[7]
port 38 nsew signal output
rlabel metal2 s 47214 99200 47270 100000 6 io_wbs_data_o[8]
port 39 nsew signal output
rlabel metal3 s 99200 52096 100000 52216 6 io_wbs_data_o[9]
port 40 nsew signal output
rlabel metal3 s 99200 11160 100000 11280 6 io_wbs_m2s_addr[0]
port 41 nsew signal input
rlabel metal3 s 99200 56584 100000 56704 6 io_wbs_m2s_addr[10]
port 42 nsew signal input
rlabel metal3 s 0 35096 800 35216 6 io_wbs_m2s_addr[11]
port 43 nsew signal input
rlabel metal2 s 63866 99200 63922 100000 6 io_wbs_m2s_addr[12]
port 44 nsew signal input
rlabel metal3 s 99200 61208 100000 61328 6 io_wbs_m2s_addr[13]
port 45 nsew signal input
rlabel metal2 s 73158 0 73214 800 6 io_wbs_m2s_addr[14]
port 46 nsew signal input
rlabel metal2 s 69386 99200 69442 100000 6 io_wbs_m2s_addr[15]
port 47 nsew signal input
rlabel metal3 s 99200 20272 100000 20392 6 io_wbs_m2s_addr[1]
port 48 nsew signal input
rlabel metal3 s 99200 33872 100000 33992 6 io_wbs_m2s_addr[2]
port 49 nsew signal input
rlabel metal3 s 99200 38496 100000 38616 6 io_wbs_m2s_addr[3]
port 50 nsew signal input
rlabel metal2 s 30470 99200 30526 100000 6 io_wbs_m2s_addr[4]
port 51 nsew signal input
rlabel metal2 s 36082 99200 36138 100000 6 io_wbs_m2s_addr[5]
port 52 nsew signal input
rlabel metal2 s 30286 0 30342 800 6 io_wbs_m2s_addr[6]
port 53 nsew signal input
rlabel metal2 s 37462 0 37518 800 6 io_wbs_m2s_addr[7]
port 54 nsew signal input
rlabel metal2 s 52734 99200 52790 100000 6 io_wbs_m2s_addr[8]
port 55 nsew signal input
rlabel metal3 s 0 31288 800 31408 6 io_wbs_m2s_addr[9]
port 56 nsew signal input
rlabel metal3 s 99200 15784 100000 15904 6 io_wbs_m2s_data[0]
port 57 nsew signal input
rlabel metal2 s 51722 0 51778 800 6 io_wbs_m2s_data[10]
port 58 nsew signal input
rlabel metal2 s 58898 0 58954 800 6 io_wbs_m2s_data[11]
port 59 nsew signal input
rlabel metal2 s 62394 0 62450 800 6 io_wbs_m2s_data[12]
port 60 nsew signal input
rlabel metal2 s 69570 0 69626 800 6 io_wbs_m2s_data[13]
port 61 nsew signal input
rlabel metal3 s 99200 70320 100000 70440 6 io_wbs_m2s_data[14]
port 62 nsew signal input
rlabel metal3 s 0 42440 800 42560 6 io_wbs_m2s_data[15]
port 63 nsew signal input
rlabel metal2 s 80334 0 80390 800 6 io_wbs_m2s_data[16]
port 64 nsew signal input
rlabel metal3 s 0 49784 800 49904 6 io_wbs_m2s_data[17]
port 65 nsew signal input
rlabel metal2 s 74998 99200 75054 100000 6 io_wbs_m2s_data[18]
port 66 nsew signal input
rlabel metal2 s 87418 0 87474 800 6 io_wbs_m2s_data[19]
port 67 nsew signal input
rlabel metal3 s 99200 24896 100000 25016 6 io_wbs_m2s_data[1]
port 68 nsew signal input
rlabel metal3 s 0 57264 800 57384 6 io_wbs_m2s_data[20]
port 69 nsew signal input
rlabel metal3 s 0 64608 800 64728 6 io_wbs_m2s_data[21]
port 70 nsew signal input
rlabel metal3 s 0 68416 800 68536 6 io_wbs_m2s_data[22]
port 71 nsew signal input
rlabel metal3 s 99200 88408 100000 88528 6 io_wbs_m2s_data[23]
port 72 nsew signal input
rlabel metal2 s 86038 99200 86094 100000 6 io_wbs_m2s_data[24]
port 73 nsew signal input
rlabel metal2 s 91650 99200 91706 100000 6 io_wbs_m2s_data[25]
port 74 nsew signal input
rlabel metal3 s 0 75760 800 75880 6 io_wbs_m2s_data[26]
port 75 nsew signal input
rlabel metal3 s 0 83104 800 83224 6 io_wbs_m2s_data[27]
port 76 nsew signal input
rlabel metal3 s 0 90584 800 90704 6 io_wbs_m2s_data[28]
port 77 nsew signal input
rlabel metal2 s 98182 0 98238 800 6 io_wbs_m2s_data[29]
port 78 nsew signal input
rlabel metal3 s 0 20272 800 20392 6 io_wbs_m2s_data[2]
port 79 nsew signal input
rlabel metal3 s 99200 97520 100000 97640 6 io_wbs_m2s_data[30]
port 80 nsew signal input
rlabel metal3 s 0 97928 800 98048 6 io_wbs_m2s_data[31]
port 81 nsew signal input
rlabel metal2 s 24950 99200 25006 100000 6 io_wbs_m2s_data[3]
port 82 nsew signal input
rlabel metal2 s 26698 0 26754 800 6 io_wbs_m2s_data[4]
port 83 nsew signal input
rlabel metal2 s 41602 99200 41658 100000 6 io_wbs_m2s_data[5]
port 84 nsew signal input
rlabel metal2 s 33874 0 33930 800 6 io_wbs_m2s_data[6]
port 85 nsew signal input
rlabel metal2 s 41050 0 41106 800 6 io_wbs_m2s_data[7]
port 86 nsew signal input
rlabel metal2 s 44546 0 44602 800 6 io_wbs_m2s_data[8]
port 87 nsew signal input
rlabel metal2 s 48134 0 48190 800 6 io_wbs_m2s_data[9]
port 88 nsew signal input
rlabel metal2 s 19430 99200 19486 100000 6 io_wbs_m2s_sel[0]
port 89 nsew signal input
rlabel metal3 s 0 16464 800 16584 6 io_wbs_m2s_sel[1]
port 90 nsew signal input
rlabel metal2 s 16026 0 16082 800 6 io_wbs_m2s_sel[2]
port 91 nsew signal input
rlabel metal3 s 0 23944 800 24064 6 io_wbs_m2s_sel[3]
port 92 nsew signal input
rlabel metal2 s 12438 0 12494 800 6 io_wbs_m2s_stb
port 93 nsew signal input
rlabel metal3 s 0 9120 800 9240 6 io_wbs_m2s_we
port 94 nsew signal input
rlabel metal2 s 5262 0 5318 800 6 reset
port 95 nsew signal input
rlabel metal4 s 4208 2128 4528 97424 6 vccd1
port 96 nsew power input
rlabel metal4 s 34928 2128 35248 97424 6 vccd1
port 96 nsew power input
rlabel metal4 s 65648 2128 65968 97424 6 vccd1
port 96 nsew power input
rlabel metal4 s 96368 2128 96688 97424 6 vccd1
port 96 nsew power input
rlabel metal4 s 19568 2128 19888 97424 6 vssd1
port 97 nsew ground input
rlabel metal4 s 50288 2128 50608 97424 6 vssd1
port 97 nsew ground input
rlabel metal4 s 81008 2128 81328 97424 6 vssd1
port 97 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 100000 100000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 17551748
string GDS_FILE /home/em/mpw/UETRV-ECORE/openlane/Motor_Top/runs/Motor_Top/results/finishing/Motor_Top.magic.gds
string GDS_START 1058546
<< end >>

