magic
tech sky130A
magscale 1 2
timestamp 1647906485
<< obsli1 >>
rect 1104 2159 98808 97393
<< obsm1 >>
rect 1104 2128 98808 97424
<< metal2 >>
rect 4986 99200 5042 100000
rect 14922 99200 14978 100000
rect 24950 99200 25006 100000
rect 34978 99200 35034 100000
rect 44914 99200 44970 100000
rect 54942 99200 54998 100000
rect 64970 99200 65026 100000
rect 74906 99200 74962 100000
rect 84934 99200 84990 100000
rect 94962 99200 95018 100000
rect 4158 0 4214 800
rect 12438 0 12494 800
rect 20810 0 20866 800
rect 29090 0 29146 800
rect 37462 0 37518 800
rect 45742 0 45798 800
rect 54114 0 54170 800
rect 62486 0 62542 800
rect 70766 0 70822 800
rect 79138 0 79194 800
rect 87418 0 87474 800
rect 95790 0 95846 800
<< obsm2 >>
rect 1398 99144 4930 99362
rect 5098 99144 14866 99362
rect 15034 99144 24894 99362
rect 25062 99144 34922 99362
rect 35090 99144 44858 99362
rect 45026 99144 54886 99362
rect 55054 99144 64914 99362
rect 65082 99144 74850 99362
rect 75018 99144 84878 99362
rect 85046 99144 94906 99362
rect 95074 99144 98238 99362
rect 1398 856 98238 99144
rect 1398 711 4102 856
rect 4270 711 12382 856
rect 12550 711 20754 856
rect 20922 711 29034 856
rect 29202 711 37406 856
rect 37574 711 45686 856
rect 45854 711 54058 856
rect 54226 711 62430 856
rect 62598 711 70710 856
rect 70878 711 79082 856
rect 79250 711 87362 856
rect 87530 711 95734 856
rect 95902 711 98238 856
<< metal3 >>
rect 0 99016 800 99136
rect 0 97520 800 97640
rect 0 95888 800 96008
rect 99200 95344 100000 95464
rect 0 94392 800 94512
rect 0 92760 800 92880
rect 0 91264 800 91384
rect 0 89632 800 89752
rect 0 88136 800 88256
rect 0 86504 800 86624
rect 99200 86232 100000 86352
rect 0 85008 800 85128
rect 0 83376 800 83496
rect 0 81880 800 82000
rect 0 80248 800 80368
rect 0 78752 800 78872
rect 0 77120 800 77240
rect 99200 77120 100000 77240
rect 0 75624 800 75744
rect 0 73992 800 74112
rect 0 72496 800 72616
rect 0 70864 800 70984
rect 0 69368 800 69488
rect 99200 68008 100000 68128
rect 0 67736 800 67856
rect 0 66240 800 66360
rect 0 64608 800 64728
rect 0 63112 800 63232
rect 0 61480 800 61600
rect 0 59984 800 60104
rect 99200 58896 100000 59016
rect 0 58352 800 58472
rect 0 56856 800 56976
rect 0 55224 800 55344
rect 0 53728 800 53848
rect 0 52096 800 52216
rect 0 50600 800 50720
rect 99200 49920 100000 50040
rect 0 49104 800 49224
rect 0 47472 800 47592
rect 0 45976 800 46096
rect 0 44344 800 44464
rect 0 42848 800 42968
rect 0 41216 800 41336
rect 99200 40808 100000 40928
rect 0 39720 800 39840
rect 0 38088 800 38208
rect 0 36592 800 36712
rect 0 34960 800 35080
rect 0 33464 800 33584
rect 0 31832 800 31952
rect 99200 31696 100000 31816
rect 0 30336 800 30456
rect 0 28704 800 28824
rect 0 27208 800 27328
rect 0 25576 800 25696
rect 0 24080 800 24200
rect 0 22448 800 22568
rect 99200 22584 100000 22704
rect 0 20952 800 21072
rect 0 19320 800 19440
rect 0 17824 800 17944
rect 0 16192 800 16312
rect 0 14696 800 14816
rect 99200 13472 100000 13592
rect 0 13064 800 13184
rect 0 11568 800 11688
rect 0 9936 800 10056
rect 0 8440 800 8560
rect 0 6808 800 6928
rect 0 5312 800 5432
rect 99200 4496 100000 4616
rect 0 3680 800 3800
rect 0 2184 800 2304
rect 0 688 800 808
<< obsm3 >>
rect 880 98936 99200 99109
rect 800 97720 99200 98936
rect 880 97440 99200 97720
rect 800 96088 99200 97440
rect 880 95808 99200 96088
rect 800 95544 99200 95808
rect 800 95264 99120 95544
rect 800 94592 99200 95264
rect 880 94312 99200 94592
rect 800 92960 99200 94312
rect 880 92680 99200 92960
rect 800 91464 99200 92680
rect 880 91184 99200 91464
rect 800 89832 99200 91184
rect 880 89552 99200 89832
rect 800 88336 99200 89552
rect 880 88056 99200 88336
rect 800 86704 99200 88056
rect 880 86432 99200 86704
rect 880 86424 99120 86432
rect 800 86152 99120 86424
rect 800 85208 99200 86152
rect 880 84928 99200 85208
rect 800 83576 99200 84928
rect 880 83296 99200 83576
rect 800 82080 99200 83296
rect 880 81800 99200 82080
rect 800 80448 99200 81800
rect 880 80168 99200 80448
rect 800 78952 99200 80168
rect 880 78672 99200 78952
rect 800 77320 99200 78672
rect 880 77040 99120 77320
rect 800 75824 99200 77040
rect 880 75544 99200 75824
rect 800 74192 99200 75544
rect 880 73912 99200 74192
rect 800 72696 99200 73912
rect 880 72416 99200 72696
rect 800 71064 99200 72416
rect 880 70784 99200 71064
rect 800 69568 99200 70784
rect 880 69288 99200 69568
rect 800 68208 99200 69288
rect 800 67936 99120 68208
rect 880 67928 99120 67936
rect 880 67656 99200 67928
rect 800 66440 99200 67656
rect 880 66160 99200 66440
rect 800 64808 99200 66160
rect 880 64528 99200 64808
rect 800 63312 99200 64528
rect 880 63032 99200 63312
rect 800 61680 99200 63032
rect 880 61400 99200 61680
rect 800 60184 99200 61400
rect 880 59904 99200 60184
rect 800 59096 99200 59904
rect 800 58816 99120 59096
rect 800 58552 99200 58816
rect 880 58272 99200 58552
rect 800 57056 99200 58272
rect 880 56776 99200 57056
rect 800 55424 99200 56776
rect 880 55144 99200 55424
rect 800 53928 99200 55144
rect 880 53648 99200 53928
rect 800 52296 99200 53648
rect 880 52016 99200 52296
rect 800 50800 99200 52016
rect 880 50520 99200 50800
rect 800 50120 99200 50520
rect 800 49840 99120 50120
rect 800 49304 99200 49840
rect 880 49024 99200 49304
rect 800 47672 99200 49024
rect 880 47392 99200 47672
rect 800 46176 99200 47392
rect 880 45896 99200 46176
rect 800 44544 99200 45896
rect 880 44264 99200 44544
rect 800 43048 99200 44264
rect 880 42768 99200 43048
rect 800 41416 99200 42768
rect 880 41136 99200 41416
rect 800 41008 99200 41136
rect 800 40728 99120 41008
rect 800 39920 99200 40728
rect 880 39640 99200 39920
rect 800 38288 99200 39640
rect 880 38008 99200 38288
rect 800 36792 99200 38008
rect 880 36512 99200 36792
rect 800 35160 99200 36512
rect 880 34880 99200 35160
rect 800 33664 99200 34880
rect 880 33384 99200 33664
rect 800 32032 99200 33384
rect 880 31896 99200 32032
rect 880 31752 99120 31896
rect 800 31616 99120 31752
rect 800 30536 99200 31616
rect 880 30256 99200 30536
rect 800 28904 99200 30256
rect 880 28624 99200 28904
rect 800 27408 99200 28624
rect 880 27128 99200 27408
rect 800 25776 99200 27128
rect 880 25496 99200 25776
rect 800 24280 99200 25496
rect 880 24000 99200 24280
rect 800 22784 99200 24000
rect 800 22648 99120 22784
rect 880 22504 99120 22648
rect 880 22368 99200 22504
rect 800 21152 99200 22368
rect 880 20872 99200 21152
rect 800 19520 99200 20872
rect 880 19240 99200 19520
rect 800 18024 99200 19240
rect 880 17744 99200 18024
rect 800 16392 99200 17744
rect 880 16112 99200 16392
rect 800 14896 99200 16112
rect 880 14616 99200 14896
rect 800 13672 99200 14616
rect 800 13392 99120 13672
rect 800 13264 99200 13392
rect 880 12984 99200 13264
rect 800 11768 99200 12984
rect 880 11488 99200 11768
rect 800 10136 99200 11488
rect 880 9856 99200 10136
rect 800 8640 99200 9856
rect 880 8360 99200 8640
rect 800 7008 99200 8360
rect 880 6728 99200 7008
rect 800 5512 99200 6728
rect 880 5232 99200 5512
rect 800 4696 99200 5232
rect 800 4416 99120 4696
rect 800 3880 99200 4416
rect 880 3600 99200 3880
rect 800 2384 99200 3600
rect 880 2104 99200 2384
rect 800 888 99200 2104
rect 880 715 99200 888
<< metal4 >>
rect 4208 2128 4528 97424
rect 19568 2128 19888 97424
rect 34928 2128 35248 97424
rect 50288 2128 50608 97424
rect 65648 2128 65968 97424
rect 81008 2128 81328 97424
rect 96368 2128 96688 97424
<< obsm4 >>
rect 8155 2619 19488 95845
rect 19968 2619 34848 95845
rect 35328 2619 50208 95845
rect 50688 2619 57901 95845
<< labels >>
rlabel metal2 s 4986 99200 5042 100000 6 clock
port 1 nsew signal input
rlabel metal3 s 0 85008 800 85128 6 io_ba_match
port 2 nsew signal input
rlabel metal2 s 20810 0 20866 800 6 io_motor_irq
port 3 nsew signal output
rlabel metal3 s 99200 4496 100000 4616 6 io_pwm_high
port 4 nsew signal output
rlabel metal3 s 99200 22584 100000 22704 6 io_pwm_high_en
port 5 nsew signal output
rlabel metal3 s 99200 13472 100000 13592 6 io_pwm_low
port 6 nsew signal output
rlabel metal2 s 24950 99200 25006 100000 6 io_pwm_low_en
port 7 nsew signal output
rlabel metal2 s 4158 0 4214 800 6 io_qei_ch_a
port 8 nsew signal input
rlabel metal2 s 12438 0 12494 800 6 io_qei_ch_b
port 9 nsew signal input
rlabel metal3 s 99200 31696 100000 31816 6 io_wbs_ack_o
port 10 nsew signal output
rlabel metal2 s 34978 99200 35034 100000 6 io_wbs_data_o[0]
port 11 nsew signal output
rlabel metal2 s 45742 0 45798 800 6 io_wbs_data_o[10]
port 12 nsew signal output
rlabel metal3 s 99200 68008 100000 68128 6 io_wbs_data_o[11]
port 13 nsew signal output
rlabel metal2 s 54114 0 54170 800 6 io_wbs_data_o[12]
port 14 nsew signal output
rlabel metal2 s 62486 0 62542 800 6 io_wbs_data_o[13]
port 15 nsew signal output
rlabel metal3 s 0 88136 800 88256 6 io_wbs_data_o[14]
port 16 nsew signal output
rlabel metal2 s 74906 99200 74962 100000 6 io_wbs_data_o[15]
port 17 nsew signal output
rlabel metal2 s 70766 0 70822 800 6 io_wbs_data_o[16]
port 18 nsew signal output
rlabel metal3 s 0 89632 800 89752 6 io_wbs_data_o[17]
port 19 nsew signal output
rlabel metal2 s 79138 0 79194 800 6 io_wbs_data_o[18]
port 20 nsew signal output
rlabel metal3 s 0 91264 800 91384 6 io_wbs_data_o[19]
port 21 nsew signal output
rlabel metal3 s 0 86504 800 86624 6 io_wbs_data_o[1]
port 22 nsew signal output
rlabel metal3 s 0 92760 800 92880 6 io_wbs_data_o[20]
port 23 nsew signal output
rlabel metal2 s 84934 99200 84990 100000 6 io_wbs_data_o[21]
port 24 nsew signal output
rlabel metal3 s 0 94392 800 94512 6 io_wbs_data_o[22]
port 25 nsew signal output
rlabel metal3 s 99200 77120 100000 77240 6 io_wbs_data_o[23]
port 26 nsew signal output
rlabel metal2 s 87418 0 87474 800 6 io_wbs_data_o[24]
port 27 nsew signal output
rlabel metal3 s 0 95888 800 96008 6 io_wbs_data_o[25]
port 28 nsew signal output
rlabel metal3 s 0 97520 800 97640 6 io_wbs_data_o[26]
port 29 nsew signal output
rlabel metal3 s 0 99016 800 99136 6 io_wbs_data_o[27]
port 30 nsew signal output
rlabel metal2 s 95790 0 95846 800 6 io_wbs_data_o[28]
port 31 nsew signal output
rlabel metal2 s 94962 99200 95018 100000 6 io_wbs_data_o[29]
port 32 nsew signal output
rlabel metal2 s 44914 99200 44970 100000 6 io_wbs_data_o[2]
port 33 nsew signal output
rlabel metal3 s 99200 86232 100000 86352 6 io_wbs_data_o[30]
port 34 nsew signal output
rlabel metal3 s 99200 95344 100000 95464 6 io_wbs_data_o[31]
port 35 nsew signal output
rlabel metal2 s 54942 99200 54998 100000 6 io_wbs_data_o[3]
port 36 nsew signal output
rlabel metal2 s 64970 99200 65026 100000 6 io_wbs_data_o[4]
port 37 nsew signal output
rlabel metal3 s 99200 40808 100000 40928 6 io_wbs_data_o[5]
port 38 nsew signal output
rlabel metal3 s 99200 49920 100000 50040 6 io_wbs_data_o[6]
port 39 nsew signal output
rlabel metal2 s 29090 0 29146 800 6 io_wbs_data_o[7]
port 40 nsew signal output
rlabel metal3 s 99200 58896 100000 59016 6 io_wbs_data_o[8]
port 41 nsew signal output
rlabel metal2 s 37462 0 37518 800 6 io_wbs_data_o[9]
port 42 nsew signal output
rlabel metal3 s 0 3680 800 3800 6 io_wbs_m2s_addr[0]
port 43 nsew signal input
rlabel metal3 s 0 41216 800 41336 6 io_wbs_m2s_addr[10]
port 44 nsew signal input
rlabel metal3 s 0 44344 800 44464 6 io_wbs_m2s_addr[11]
port 45 nsew signal input
rlabel metal3 s 0 47472 800 47592 6 io_wbs_m2s_addr[12]
port 46 nsew signal input
rlabel metal3 s 0 50600 800 50720 6 io_wbs_m2s_addr[13]
port 47 nsew signal input
rlabel metal3 s 0 53728 800 53848 6 io_wbs_m2s_addr[14]
port 48 nsew signal input
rlabel metal3 s 0 56856 800 56976 6 io_wbs_m2s_addr[15]
port 49 nsew signal input
rlabel metal3 s 0 8440 800 8560 6 io_wbs_m2s_addr[1]
port 50 nsew signal input
rlabel metal3 s 0 13064 800 13184 6 io_wbs_m2s_addr[2]
port 51 nsew signal input
rlabel metal3 s 0 17824 800 17944 6 io_wbs_m2s_addr[3]
port 52 nsew signal input
rlabel metal3 s 0 22448 800 22568 6 io_wbs_m2s_addr[4]
port 53 nsew signal input
rlabel metal3 s 0 25576 800 25696 6 io_wbs_m2s_addr[5]
port 54 nsew signal input
rlabel metal3 s 0 28704 800 28824 6 io_wbs_m2s_addr[6]
port 55 nsew signal input
rlabel metal3 s 0 31832 800 31952 6 io_wbs_m2s_addr[7]
port 56 nsew signal input
rlabel metal3 s 0 34960 800 35080 6 io_wbs_m2s_addr[8]
port 57 nsew signal input
rlabel metal3 s 0 38088 800 38208 6 io_wbs_m2s_addr[9]
port 58 nsew signal input
rlabel metal3 s 0 5312 800 5432 6 io_wbs_m2s_data[0]
port 59 nsew signal input
rlabel metal3 s 0 42848 800 42968 6 io_wbs_m2s_data[10]
port 60 nsew signal input
rlabel metal3 s 0 45976 800 46096 6 io_wbs_m2s_data[11]
port 61 nsew signal input
rlabel metal3 s 0 49104 800 49224 6 io_wbs_m2s_data[12]
port 62 nsew signal input
rlabel metal3 s 0 52096 800 52216 6 io_wbs_m2s_data[13]
port 63 nsew signal input
rlabel metal3 s 0 55224 800 55344 6 io_wbs_m2s_data[14]
port 64 nsew signal input
rlabel metal3 s 0 58352 800 58472 6 io_wbs_m2s_data[15]
port 65 nsew signal input
rlabel metal3 s 0 59984 800 60104 6 io_wbs_m2s_data[16]
port 66 nsew signal input
rlabel metal3 s 0 61480 800 61600 6 io_wbs_m2s_data[17]
port 67 nsew signal input
rlabel metal3 s 0 63112 800 63232 6 io_wbs_m2s_data[18]
port 68 nsew signal input
rlabel metal3 s 0 64608 800 64728 6 io_wbs_m2s_data[19]
port 69 nsew signal input
rlabel metal3 s 0 9936 800 10056 6 io_wbs_m2s_data[1]
port 70 nsew signal input
rlabel metal3 s 0 66240 800 66360 6 io_wbs_m2s_data[20]
port 71 nsew signal input
rlabel metal3 s 0 67736 800 67856 6 io_wbs_m2s_data[21]
port 72 nsew signal input
rlabel metal3 s 0 69368 800 69488 6 io_wbs_m2s_data[22]
port 73 nsew signal input
rlabel metal3 s 0 70864 800 70984 6 io_wbs_m2s_data[23]
port 74 nsew signal input
rlabel metal3 s 0 72496 800 72616 6 io_wbs_m2s_data[24]
port 75 nsew signal input
rlabel metal3 s 0 73992 800 74112 6 io_wbs_m2s_data[25]
port 76 nsew signal input
rlabel metal3 s 0 75624 800 75744 6 io_wbs_m2s_data[26]
port 77 nsew signal input
rlabel metal3 s 0 77120 800 77240 6 io_wbs_m2s_data[27]
port 78 nsew signal input
rlabel metal3 s 0 78752 800 78872 6 io_wbs_m2s_data[28]
port 79 nsew signal input
rlabel metal3 s 0 80248 800 80368 6 io_wbs_m2s_data[29]
port 80 nsew signal input
rlabel metal3 s 0 14696 800 14816 6 io_wbs_m2s_data[2]
port 81 nsew signal input
rlabel metal3 s 0 81880 800 82000 6 io_wbs_m2s_data[30]
port 82 nsew signal input
rlabel metal3 s 0 83376 800 83496 6 io_wbs_m2s_data[31]
port 83 nsew signal input
rlabel metal3 s 0 19320 800 19440 6 io_wbs_m2s_data[3]
port 84 nsew signal input
rlabel metal3 s 0 24080 800 24200 6 io_wbs_m2s_data[4]
port 85 nsew signal input
rlabel metal3 s 0 27208 800 27328 6 io_wbs_m2s_data[5]
port 86 nsew signal input
rlabel metal3 s 0 30336 800 30456 6 io_wbs_m2s_data[6]
port 87 nsew signal input
rlabel metal3 s 0 33464 800 33584 6 io_wbs_m2s_data[7]
port 88 nsew signal input
rlabel metal3 s 0 36592 800 36712 6 io_wbs_m2s_data[8]
port 89 nsew signal input
rlabel metal3 s 0 39720 800 39840 6 io_wbs_m2s_data[9]
port 90 nsew signal input
rlabel metal3 s 0 6808 800 6928 6 io_wbs_m2s_sel[0]
port 91 nsew signal input
rlabel metal3 s 0 11568 800 11688 6 io_wbs_m2s_sel[1]
port 92 nsew signal input
rlabel metal3 s 0 16192 800 16312 6 io_wbs_m2s_sel[2]
port 93 nsew signal input
rlabel metal3 s 0 20952 800 21072 6 io_wbs_m2s_sel[3]
port 94 nsew signal input
rlabel metal3 s 0 688 800 808 6 io_wbs_m2s_stb
port 95 nsew signal input
rlabel metal3 s 0 2184 800 2304 6 io_wbs_m2s_we
port 96 nsew signal input
rlabel metal2 s 14922 99200 14978 100000 6 reset
port 97 nsew signal input
rlabel metal4 s 4208 2128 4528 97424 6 vccd1
port 98 nsew power input
rlabel metal4 s 34928 2128 35248 97424 6 vccd1
port 98 nsew power input
rlabel metal4 s 65648 2128 65968 97424 6 vccd1
port 98 nsew power input
rlabel metal4 s 96368 2128 96688 97424 6 vccd1
port 98 nsew power input
rlabel metal4 s 19568 2128 19888 97424 6 vssd1
port 99 nsew ground input
rlabel metal4 s 50288 2128 50608 97424 6 vssd1
port 99 nsew ground input
rlabel metal4 s 81008 2128 81328 97424 6 vssd1
port 99 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 100000 100000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 17666050
string GDS_FILE /home/ali112000/mpw5/UETRV-ECORE/openlane/Motor_Top/runs/Motor_Top/results/finishing/Motor_Top.magic.gds
string GDS_START 1110772
<< end >>

