magic
tech sky130A
magscale 1 2
timestamp 1649143826
<< obsli1 >>
rect 1104 2159 218868 217617
<< obsm1 >>
rect 1104 1980 219130 217648
<< metal2 >>
rect 846 219200 902 220000
rect 2502 219200 2558 220000
rect 4250 219200 4306 220000
rect 5998 219200 6054 220000
rect 7746 219200 7802 220000
rect 9494 219200 9550 220000
rect 11242 219200 11298 220000
rect 12990 219200 13046 220000
rect 14738 219200 14794 220000
rect 16486 219200 16542 220000
rect 18234 219200 18290 220000
rect 19982 219200 20038 220000
rect 21730 219200 21786 220000
rect 23478 219200 23534 220000
rect 25226 219200 25282 220000
rect 26974 219200 27030 220000
rect 28722 219200 28778 220000
rect 30470 219200 30526 220000
rect 32218 219200 32274 220000
rect 33966 219200 34022 220000
rect 35714 219200 35770 220000
rect 37462 219200 37518 220000
rect 39210 219200 39266 220000
rect 40958 219200 41014 220000
rect 42706 219200 42762 220000
rect 44454 219200 44510 220000
rect 46202 219200 46258 220000
rect 47950 219200 48006 220000
rect 49698 219200 49754 220000
rect 51446 219200 51502 220000
rect 53194 219200 53250 220000
rect 54942 219200 54998 220000
rect 56690 219200 56746 220000
rect 58438 219200 58494 220000
rect 60186 219200 60242 220000
rect 61934 219200 61990 220000
rect 63682 219200 63738 220000
rect 65430 219200 65486 220000
rect 67178 219200 67234 220000
rect 68926 219200 68982 220000
rect 70674 219200 70730 220000
rect 72422 219200 72478 220000
rect 74170 219200 74226 220000
rect 75826 219200 75882 220000
rect 77574 219200 77630 220000
rect 79322 219200 79378 220000
rect 81070 219200 81126 220000
rect 82818 219200 82874 220000
rect 84566 219200 84622 220000
rect 86314 219200 86370 220000
rect 88062 219200 88118 220000
rect 89810 219200 89866 220000
rect 91558 219200 91614 220000
rect 93306 219200 93362 220000
rect 95054 219200 95110 220000
rect 96802 219200 96858 220000
rect 98550 219200 98606 220000
rect 100298 219200 100354 220000
rect 102046 219200 102102 220000
rect 103794 219200 103850 220000
rect 105542 219200 105598 220000
rect 107290 219200 107346 220000
rect 109038 219200 109094 220000
rect 110786 219200 110842 220000
rect 112534 219200 112590 220000
rect 114282 219200 114338 220000
rect 116030 219200 116086 220000
rect 117778 219200 117834 220000
rect 119526 219200 119582 220000
rect 121274 219200 121330 220000
rect 123022 219200 123078 220000
rect 124770 219200 124826 220000
rect 126518 219200 126574 220000
rect 128266 219200 128322 220000
rect 130014 219200 130070 220000
rect 131762 219200 131818 220000
rect 133510 219200 133566 220000
rect 135258 219200 135314 220000
rect 137006 219200 137062 220000
rect 138754 219200 138810 220000
rect 140502 219200 140558 220000
rect 142250 219200 142306 220000
rect 143998 219200 144054 220000
rect 145746 219200 145802 220000
rect 147494 219200 147550 220000
rect 149150 219200 149206 220000
rect 150898 219200 150954 220000
rect 152646 219200 152702 220000
rect 154394 219200 154450 220000
rect 156142 219200 156198 220000
rect 157890 219200 157946 220000
rect 159638 219200 159694 220000
rect 161386 219200 161442 220000
rect 163134 219200 163190 220000
rect 164882 219200 164938 220000
rect 166630 219200 166686 220000
rect 168378 219200 168434 220000
rect 170126 219200 170182 220000
rect 171874 219200 171930 220000
rect 173622 219200 173678 220000
rect 175370 219200 175426 220000
rect 177118 219200 177174 220000
rect 178866 219200 178922 220000
rect 180614 219200 180670 220000
rect 182362 219200 182418 220000
rect 184110 219200 184166 220000
rect 185858 219200 185914 220000
rect 187606 219200 187662 220000
rect 189354 219200 189410 220000
rect 191102 219200 191158 220000
rect 192850 219200 192906 220000
rect 194598 219200 194654 220000
rect 196346 219200 196402 220000
rect 198094 219200 198150 220000
rect 199842 219200 199898 220000
rect 201590 219200 201646 220000
rect 203338 219200 203394 220000
rect 205086 219200 205142 220000
rect 206834 219200 206890 220000
rect 208582 219200 208638 220000
rect 210330 219200 210386 220000
rect 212078 219200 212134 220000
rect 213826 219200 213882 220000
rect 215574 219200 215630 220000
rect 217322 219200 217378 220000
rect 219070 219200 219126 220000
rect 1950 0 2006 800
rect 5906 0 5962 800
rect 9862 0 9918 800
rect 13910 0 13966 800
rect 17866 0 17922 800
rect 21914 0 21970 800
rect 25870 0 25926 800
rect 29918 0 29974 800
rect 33874 0 33930 800
rect 37922 0 37978 800
rect 41878 0 41934 800
rect 45926 0 45982 800
rect 49882 0 49938 800
rect 53930 0 53986 800
rect 57886 0 57942 800
rect 61934 0 61990 800
rect 65890 0 65946 800
rect 69938 0 69994 800
rect 73894 0 73950 800
rect 77850 0 77906 800
rect 81898 0 81954 800
rect 85854 0 85910 800
rect 89902 0 89958 800
rect 93858 0 93914 800
rect 97906 0 97962 800
rect 101862 0 101918 800
rect 105910 0 105966 800
rect 109866 0 109922 800
rect 113914 0 113970 800
rect 117870 0 117926 800
rect 121918 0 121974 800
rect 125874 0 125930 800
rect 129922 0 129978 800
rect 133878 0 133934 800
rect 137926 0 137982 800
rect 141882 0 141938 800
rect 145930 0 145986 800
rect 149886 0 149942 800
rect 153842 0 153898 800
rect 157890 0 157946 800
rect 161846 0 161902 800
rect 165894 0 165950 800
rect 169850 0 169906 800
rect 173898 0 173954 800
rect 177854 0 177910 800
rect 181902 0 181958 800
rect 185858 0 185914 800
rect 189906 0 189962 800
rect 193862 0 193918 800
rect 197910 0 197966 800
rect 201866 0 201922 800
rect 205914 0 205970 800
rect 209870 0 209926 800
rect 213918 0 213974 800
rect 217874 0 217930 800
<< obsm2 >>
rect 958 219144 2446 219473
rect 2614 219144 4194 219473
rect 4362 219144 5942 219473
rect 6110 219144 7690 219473
rect 7858 219144 9438 219473
rect 9606 219144 11186 219473
rect 11354 219144 12934 219473
rect 13102 219144 14682 219473
rect 14850 219144 16430 219473
rect 16598 219144 18178 219473
rect 18346 219144 19926 219473
rect 20094 219144 21674 219473
rect 21842 219144 23422 219473
rect 23590 219144 25170 219473
rect 25338 219144 26918 219473
rect 27086 219144 28666 219473
rect 28834 219144 30414 219473
rect 30582 219144 32162 219473
rect 32330 219144 33910 219473
rect 34078 219144 35658 219473
rect 35826 219144 37406 219473
rect 37574 219144 39154 219473
rect 39322 219144 40902 219473
rect 41070 219144 42650 219473
rect 42818 219144 44398 219473
rect 44566 219144 46146 219473
rect 46314 219144 47894 219473
rect 48062 219144 49642 219473
rect 49810 219144 51390 219473
rect 51558 219144 53138 219473
rect 53306 219144 54886 219473
rect 55054 219144 56634 219473
rect 56802 219144 58382 219473
rect 58550 219144 60130 219473
rect 60298 219144 61878 219473
rect 62046 219144 63626 219473
rect 63794 219144 65374 219473
rect 65542 219144 67122 219473
rect 67290 219144 68870 219473
rect 69038 219144 70618 219473
rect 70786 219144 72366 219473
rect 72534 219144 74114 219473
rect 74282 219144 75770 219473
rect 75938 219144 77518 219473
rect 77686 219144 79266 219473
rect 79434 219144 81014 219473
rect 81182 219144 82762 219473
rect 82930 219144 84510 219473
rect 84678 219144 86258 219473
rect 86426 219144 88006 219473
rect 88174 219144 89754 219473
rect 89922 219144 91502 219473
rect 91670 219144 93250 219473
rect 93418 219144 94998 219473
rect 95166 219144 96746 219473
rect 96914 219144 98494 219473
rect 98662 219144 100242 219473
rect 100410 219144 101990 219473
rect 102158 219144 103738 219473
rect 103906 219144 105486 219473
rect 105654 219144 107234 219473
rect 107402 219144 108982 219473
rect 109150 219144 110730 219473
rect 110898 219144 112478 219473
rect 112646 219144 114226 219473
rect 114394 219144 115974 219473
rect 116142 219144 117722 219473
rect 117890 219144 119470 219473
rect 119638 219144 121218 219473
rect 121386 219144 122966 219473
rect 123134 219144 124714 219473
rect 124882 219144 126462 219473
rect 126630 219144 128210 219473
rect 128378 219144 129958 219473
rect 130126 219144 131706 219473
rect 131874 219144 133454 219473
rect 133622 219144 135202 219473
rect 135370 219144 136950 219473
rect 137118 219144 138698 219473
rect 138866 219144 140446 219473
rect 140614 219144 142194 219473
rect 142362 219144 143942 219473
rect 144110 219144 145690 219473
rect 145858 219144 147438 219473
rect 147606 219144 149094 219473
rect 149262 219144 150842 219473
rect 151010 219144 152590 219473
rect 152758 219144 154338 219473
rect 154506 219144 156086 219473
rect 156254 219144 157834 219473
rect 158002 219144 159582 219473
rect 159750 219144 161330 219473
rect 161498 219144 163078 219473
rect 163246 219144 164826 219473
rect 164994 219144 166574 219473
rect 166742 219144 168322 219473
rect 168490 219144 170070 219473
rect 170238 219144 171818 219473
rect 171986 219144 173566 219473
rect 173734 219144 175314 219473
rect 175482 219144 177062 219473
rect 177230 219144 178810 219473
rect 178978 219144 180558 219473
rect 180726 219144 182306 219473
rect 182474 219144 184054 219473
rect 184222 219144 185802 219473
rect 185970 219144 187550 219473
rect 187718 219144 189298 219473
rect 189466 219144 191046 219473
rect 191214 219144 192794 219473
rect 192962 219144 194542 219473
rect 194710 219144 196290 219473
rect 196458 219144 198038 219473
rect 198206 219144 199786 219473
rect 199954 219144 201534 219473
rect 201702 219144 203282 219473
rect 203450 219144 205030 219473
rect 205198 219144 206778 219473
rect 206946 219144 208526 219473
rect 208694 219144 210274 219473
rect 210442 219144 212022 219473
rect 212190 219144 213770 219473
rect 213938 219144 215518 219473
rect 215686 219144 217266 219473
rect 217434 219144 219014 219473
rect 902 856 219124 219144
rect 902 439 1894 856
rect 2062 439 5850 856
rect 6018 439 9806 856
rect 9974 439 13854 856
rect 14022 439 17810 856
rect 17978 439 21858 856
rect 22026 439 25814 856
rect 25982 439 29862 856
rect 30030 439 33818 856
rect 33986 439 37866 856
rect 38034 439 41822 856
rect 41990 439 45870 856
rect 46038 439 49826 856
rect 49994 439 53874 856
rect 54042 439 57830 856
rect 57998 439 61878 856
rect 62046 439 65834 856
rect 66002 439 69882 856
rect 70050 439 73838 856
rect 74006 439 77794 856
rect 77962 439 81842 856
rect 82010 439 85798 856
rect 85966 439 89846 856
rect 90014 439 93802 856
rect 93970 439 97850 856
rect 98018 439 101806 856
rect 101974 439 105854 856
rect 106022 439 109810 856
rect 109978 439 113858 856
rect 114026 439 117814 856
rect 117982 439 121862 856
rect 122030 439 125818 856
rect 125986 439 129866 856
rect 130034 439 133822 856
rect 133990 439 137870 856
rect 138038 439 141826 856
rect 141994 439 145874 856
rect 146042 439 149830 856
rect 149998 439 153786 856
rect 153954 439 157834 856
rect 158002 439 161790 856
rect 161958 439 165838 856
rect 166006 439 169794 856
rect 169962 439 173842 856
rect 174010 439 177798 856
rect 177966 439 181846 856
rect 182014 439 185802 856
rect 185970 439 189850 856
rect 190018 439 193806 856
rect 193974 439 197854 856
rect 198022 439 201810 856
rect 201978 439 205858 856
rect 206026 439 209814 856
rect 209982 439 213862 856
rect 214030 439 217818 856
rect 217986 439 219124 856
<< metal3 >>
rect 0 219376 800 219496
rect 219200 218832 220000 218952
rect 0 218288 800 218408
rect 0 217200 800 217320
rect 219200 216792 220000 216912
rect 0 216248 800 216368
rect 0 215160 800 215280
rect 219200 214752 220000 214872
rect 0 214072 800 214192
rect 0 212984 800 213104
rect 219200 212712 220000 212832
rect 0 212032 800 212152
rect 0 210944 800 211064
rect 219200 210672 220000 210792
rect 0 209856 800 209976
rect 0 208768 800 208888
rect 219200 208632 220000 208752
rect 0 207816 800 207936
rect 0 206728 800 206848
rect 219200 206592 220000 206712
rect 0 205640 800 205760
rect 0 204552 800 204672
rect 219200 204552 220000 204672
rect 0 203600 800 203720
rect 0 202512 800 202632
rect 219200 202376 220000 202496
rect 0 201424 800 201544
rect 0 200336 800 200456
rect 219200 200336 220000 200456
rect 0 199384 800 199504
rect 0 198296 800 198416
rect 219200 198296 220000 198416
rect 0 197208 800 197328
rect 0 196120 800 196240
rect 219200 196256 220000 196376
rect 0 195168 800 195288
rect 0 194080 800 194200
rect 219200 194216 220000 194336
rect 0 192992 800 193112
rect 219200 192176 220000 192296
rect 0 191904 800 192024
rect 0 190952 800 191072
rect 219200 190136 220000 190256
rect 0 189864 800 189984
rect 0 188776 800 188896
rect 219200 188096 220000 188216
rect 0 187824 800 187944
rect 0 186736 800 186856
rect 219200 185920 220000 186040
rect 0 185648 800 185768
rect 0 184560 800 184680
rect 219200 183880 220000 184000
rect 0 183608 800 183728
rect 0 182520 800 182640
rect 219200 181840 220000 181960
rect 0 181432 800 181552
rect 0 180344 800 180464
rect 219200 179800 220000 179920
rect 0 179392 800 179512
rect 0 178304 800 178424
rect 219200 177760 220000 177880
rect 0 177216 800 177336
rect 0 176128 800 176248
rect 219200 175720 220000 175840
rect 0 175176 800 175296
rect 0 174088 800 174208
rect 219200 173680 220000 173800
rect 0 173000 800 173120
rect 0 171912 800 172032
rect 219200 171640 220000 171760
rect 0 170960 800 171080
rect 0 169872 800 169992
rect 219200 169464 220000 169584
rect 0 168784 800 168904
rect 0 167696 800 167816
rect 219200 167424 220000 167544
rect 0 166744 800 166864
rect 0 165656 800 165776
rect 219200 165384 220000 165504
rect 0 164568 800 164688
rect 0 163480 800 163600
rect 219200 163344 220000 163464
rect 0 162528 800 162648
rect 0 161440 800 161560
rect 219200 161304 220000 161424
rect 0 160352 800 160472
rect 0 159264 800 159384
rect 219200 159264 220000 159384
rect 0 158312 800 158432
rect 0 157224 800 157344
rect 219200 157224 220000 157344
rect 0 156136 800 156256
rect 0 155184 800 155304
rect 219200 155184 220000 155304
rect 0 154096 800 154216
rect 0 153008 800 153128
rect 219200 153008 220000 153128
rect 0 151920 800 152040
rect 0 150968 800 151088
rect 219200 150968 220000 151088
rect 0 149880 800 150000
rect 0 148792 800 148912
rect 219200 148928 220000 149048
rect 0 147704 800 147824
rect 0 146752 800 146872
rect 219200 146888 220000 147008
rect 0 145664 800 145784
rect 219200 144848 220000 144968
rect 0 144576 800 144696
rect 0 143488 800 143608
rect 219200 142808 220000 142928
rect 0 142536 800 142656
rect 0 141448 800 141568
rect 219200 140768 220000 140888
rect 0 140360 800 140480
rect 0 139272 800 139392
rect 219200 138728 220000 138848
rect 0 138320 800 138440
rect 0 137232 800 137352
rect 219200 136688 220000 136808
rect 0 136144 800 136264
rect 0 135056 800 135176
rect 219200 134512 220000 134632
rect 0 134104 800 134224
rect 0 133016 800 133136
rect 219200 132472 220000 132592
rect 0 131928 800 132048
rect 0 130840 800 130960
rect 219200 130432 220000 130552
rect 0 129888 800 130008
rect 0 128800 800 128920
rect 219200 128392 220000 128512
rect 0 127712 800 127832
rect 0 126624 800 126744
rect 219200 126352 220000 126472
rect 0 125672 800 125792
rect 0 124584 800 124704
rect 219200 124312 220000 124432
rect 0 123496 800 123616
rect 0 122544 800 122664
rect 219200 122272 220000 122392
rect 0 121456 800 121576
rect 0 120368 800 120488
rect 219200 120232 220000 120352
rect 0 119280 800 119400
rect 0 118328 800 118448
rect 219200 118056 220000 118176
rect 0 117240 800 117360
rect 0 116152 800 116272
rect 219200 116016 220000 116136
rect 0 115064 800 115184
rect 0 114112 800 114232
rect 219200 113976 220000 114096
rect 0 113024 800 113144
rect 0 111936 800 112056
rect 219200 111936 220000 112056
rect 0 110848 800 110968
rect 0 109896 800 110016
rect 219200 109896 220000 110016
rect 0 108808 800 108928
rect 0 107720 800 107840
rect 219200 107856 220000 107976
rect 0 106632 800 106752
rect 0 105680 800 105800
rect 219200 105816 220000 105936
rect 0 104592 800 104712
rect 219200 103776 220000 103896
rect 0 103504 800 103624
rect 0 102416 800 102536
rect 0 101464 800 101584
rect 219200 101600 220000 101720
rect 0 100376 800 100496
rect 219200 99560 220000 99680
rect 0 99288 800 99408
rect 0 98200 800 98320
rect 219200 97520 220000 97640
rect 0 97248 800 97368
rect 0 96160 800 96280
rect 219200 95480 220000 95600
rect 0 95072 800 95192
rect 0 94120 800 94240
rect 219200 93440 220000 93560
rect 0 93032 800 93152
rect 0 91944 800 92064
rect 219200 91400 220000 91520
rect 0 90856 800 90976
rect 0 89904 800 90024
rect 219200 89360 220000 89480
rect 0 88816 800 88936
rect 0 87728 800 87848
rect 219200 87320 220000 87440
rect 0 86640 800 86760
rect 0 85688 800 85808
rect 219200 85144 220000 85264
rect 0 84600 800 84720
rect 0 83512 800 83632
rect 219200 83104 220000 83224
rect 0 82424 800 82544
rect 0 81472 800 81592
rect 219200 81064 220000 81184
rect 0 80384 800 80504
rect 0 79296 800 79416
rect 219200 79024 220000 79144
rect 0 78208 800 78328
rect 0 77256 800 77376
rect 219200 76984 220000 77104
rect 0 76168 800 76288
rect 0 75080 800 75200
rect 219200 74944 220000 75064
rect 0 73992 800 74112
rect 0 73040 800 73160
rect 219200 72904 220000 73024
rect 0 71952 800 72072
rect 0 70864 800 70984
rect 219200 70864 220000 70984
rect 0 69776 800 69896
rect 0 68824 800 68944
rect 219200 68824 220000 68944
rect 0 67736 800 67856
rect 0 66648 800 66768
rect 219200 66648 220000 66768
rect 0 65560 800 65680
rect 0 64608 800 64728
rect 219200 64608 220000 64728
rect 0 63520 800 63640
rect 0 62432 800 62552
rect 219200 62568 220000 62688
rect 0 61480 800 61600
rect 0 60392 800 60512
rect 219200 60528 220000 60648
rect 0 59304 800 59424
rect 219200 58488 220000 58608
rect 0 58216 800 58336
rect 0 57264 800 57384
rect 219200 56448 220000 56568
rect 0 56176 800 56296
rect 0 55088 800 55208
rect 219200 54408 220000 54528
rect 0 54000 800 54120
rect 0 53048 800 53168
rect 219200 52368 220000 52488
rect 0 51960 800 52080
rect 0 50872 800 50992
rect 219200 50192 220000 50312
rect 0 49784 800 49904
rect 0 48832 800 48952
rect 219200 48152 220000 48272
rect 0 47744 800 47864
rect 0 46656 800 46776
rect 219200 46112 220000 46232
rect 0 45568 800 45688
rect 0 44616 800 44736
rect 219200 44072 220000 44192
rect 0 43528 800 43648
rect 0 42440 800 42560
rect 219200 42032 220000 42152
rect 0 41352 800 41472
rect 0 40400 800 40520
rect 219200 39992 220000 40112
rect 0 39312 800 39432
rect 0 38224 800 38344
rect 219200 37952 220000 38072
rect 0 37136 800 37256
rect 0 36184 800 36304
rect 219200 35912 220000 36032
rect 0 35096 800 35216
rect 0 34008 800 34128
rect 219200 33736 220000 33856
rect 0 32920 800 33040
rect 0 31968 800 32088
rect 219200 31696 220000 31816
rect 0 30880 800 31000
rect 0 29792 800 29912
rect 219200 29656 220000 29776
rect 0 28840 800 28960
rect 0 27752 800 27872
rect 219200 27616 220000 27736
rect 0 26664 800 26784
rect 0 25576 800 25696
rect 219200 25576 220000 25696
rect 0 24624 800 24744
rect 0 23536 800 23656
rect 219200 23536 220000 23656
rect 0 22448 800 22568
rect 0 21360 800 21480
rect 219200 21496 220000 21616
rect 0 20408 800 20528
rect 0 19320 800 19440
rect 219200 19456 220000 19576
rect 0 18232 800 18352
rect 0 17144 800 17264
rect 219200 17280 220000 17400
rect 0 16192 800 16312
rect 0 15104 800 15224
rect 219200 15240 220000 15360
rect 0 14016 800 14136
rect 219200 13200 220000 13320
rect 0 12928 800 13048
rect 0 11976 800 12096
rect 219200 11160 220000 11280
rect 0 10888 800 11008
rect 0 9800 800 9920
rect 219200 9120 220000 9240
rect 0 8712 800 8832
rect 0 7760 800 7880
rect 219200 7080 220000 7200
rect 0 6672 800 6792
rect 0 5584 800 5704
rect 219200 5040 220000 5160
rect 0 4496 800 4616
rect 0 3544 800 3664
rect 219200 3000 220000 3120
rect 0 2456 800 2576
rect 0 1368 800 1488
rect 219200 960 220000 1080
rect 0 416 800 536
<< obsm3 >>
rect 880 219296 219200 219469
rect 800 219032 219200 219296
rect 800 218752 219120 219032
rect 800 218488 219200 218752
rect 880 218208 219200 218488
rect 800 217400 219200 218208
rect 880 217120 219200 217400
rect 800 216992 219200 217120
rect 800 216712 219120 216992
rect 800 216448 219200 216712
rect 880 216168 219200 216448
rect 800 215360 219200 216168
rect 880 215080 219200 215360
rect 800 214952 219200 215080
rect 800 214672 219120 214952
rect 800 214272 219200 214672
rect 880 213992 219200 214272
rect 800 213184 219200 213992
rect 880 212912 219200 213184
rect 880 212904 219120 212912
rect 800 212632 219120 212904
rect 800 212232 219200 212632
rect 880 211952 219200 212232
rect 800 211144 219200 211952
rect 880 210872 219200 211144
rect 880 210864 219120 210872
rect 800 210592 219120 210864
rect 800 210056 219200 210592
rect 880 209776 219200 210056
rect 800 208968 219200 209776
rect 880 208832 219200 208968
rect 880 208688 219120 208832
rect 800 208552 219120 208688
rect 800 208016 219200 208552
rect 880 207736 219200 208016
rect 800 206928 219200 207736
rect 880 206792 219200 206928
rect 880 206648 219120 206792
rect 800 206512 219120 206648
rect 800 205840 219200 206512
rect 880 205560 219200 205840
rect 800 204752 219200 205560
rect 880 204472 219120 204752
rect 800 203800 219200 204472
rect 880 203520 219200 203800
rect 800 202712 219200 203520
rect 880 202576 219200 202712
rect 880 202432 219120 202576
rect 800 202296 219120 202432
rect 800 201624 219200 202296
rect 880 201344 219200 201624
rect 800 200536 219200 201344
rect 880 200256 219120 200536
rect 800 199584 219200 200256
rect 880 199304 219200 199584
rect 800 198496 219200 199304
rect 880 198216 219120 198496
rect 800 197408 219200 198216
rect 880 197128 219200 197408
rect 800 196456 219200 197128
rect 800 196320 219120 196456
rect 880 196176 219120 196320
rect 880 196040 219200 196176
rect 800 195368 219200 196040
rect 880 195088 219200 195368
rect 800 194416 219200 195088
rect 800 194280 219120 194416
rect 880 194136 219120 194280
rect 880 194000 219200 194136
rect 800 193192 219200 194000
rect 880 192912 219200 193192
rect 800 192376 219200 192912
rect 800 192104 219120 192376
rect 880 192096 219120 192104
rect 880 191824 219200 192096
rect 800 191152 219200 191824
rect 880 190872 219200 191152
rect 800 190336 219200 190872
rect 800 190064 219120 190336
rect 880 190056 219120 190064
rect 880 189784 219200 190056
rect 800 188976 219200 189784
rect 880 188696 219200 188976
rect 800 188296 219200 188696
rect 800 188024 219120 188296
rect 880 188016 219120 188024
rect 880 187744 219200 188016
rect 800 186936 219200 187744
rect 880 186656 219200 186936
rect 800 186120 219200 186656
rect 800 185848 219120 186120
rect 880 185840 219120 185848
rect 880 185568 219200 185840
rect 800 184760 219200 185568
rect 880 184480 219200 184760
rect 800 184080 219200 184480
rect 800 183808 219120 184080
rect 880 183800 219120 183808
rect 880 183528 219200 183800
rect 800 182720 219200 183528
rect 880 182440 219200 182720
rect 800 182040 219200 182440
rect 800 181760 219120 182040
rect 800 181632 219200 181760
rect 880 181352 219200 181632
rect 800 180544 219200 181352
rect 880 180264 219200 180544
rect 800 180000 219200 180264
rect 800 179720 219120 180000
rect 800 179592 219200 179720
rect 880 179312 219200 179592
rect 800 178504 219200 179312
rect 880 178224 219200 178504
rect 800 177960 219200 178224
rect 800 177680 219120 177960
rect 800 177416 219200 177680
rect 880 177136 219200 177416
rect 800 176328 219200 177136
rect 880 176048 219200 176328
rect 800 175920 219200 176048
rect 800 175640 219120 175920
rect 800 175376 219200 175640
rect 880 175096 219200 175376
rect 800 174288 219200 175096
rect 880 174008 219200 174288
rect 800 173880 219200 174008
rect 800 173600 219120 173880
rect 800 173200 219200 173600
rect 880 172920 219200 173200
rect 800 172112 219200 172920
rect 880 171840 219200 172112
rect 880 171832 219120 171840
rect 800 171560 219120 171832
rect 800 171160 219200 171560
rect 880 170880 219200 171160
rect 800 170072 219200 170880
rect 880 169792 219200 170072
rect 800 169664 219200 169792
rect 800 169384 219120 169664
rect 800 168984 219200 169384
rect 880 168704 219200 168984
rect 800 167896 219200 168704
rect 880 167624 219200 167896
rect 880 167616 219120 167624
rect 800 167344 219120 167616
rect 800 166944 219200 167344
rect 880 166664 219200 166944
rect 800 165856 219200 166664
rect 880 165584 219200 165856
rect 880 165576 219120 165584
rect 800 165304 219120 165576
rect 800 164768 219200 165304
rect 880 164488 219200 164768
rect 800 163680 219200 164488
rect 880 163544 219200 163680
rect 880 163400 219120 163544
rect 800 163264 219120 163400
rect 800 162728 219200 163264
rect 880 162448 219200 162728
rect 800 161640 219200 162448
rect 880 161504 219200 161640
rect 880 161360 219120 161504
rect 800 161224 219120 161360
rect 800 160552 219200 161224
rect 880 160272 219200 160552
rect 800 159464 219200 160272
rect 880 159184 219120 159464
rect 800 158512 219200 159184
rect 880 158232 219200 158512
rect 800 157424 219200 158232
rect 880 157144 219120 157424
rect 800 156336 219200 157144
rect 880 156056 219200 156336
rect 800 155384 219200 156056
rect 880 155104 219120 155384
rect 800 154296 219200 155104
rect 880 154016 219200 154296
rect 800 153208 219200 154016
rect 880 152928 219120 153208
rect 800 152120 219200 152928
rect 880 151840 219200 152120
rect 800 151168 219200 151840
rect 880 150888 219120 151168
rect 800 150080 219200 150888
rect 880 149800 219200 150080
rect 800 149128 219200 149800
rect 800 148992 219120 149128
rect 880 148848 219120 148992
rect 880 148712 219200 148848
rect 800 147904 219200 148712
rect 880 147624 219200 147904
rect 800 147088 219200 147624
rect 800 146952 219120 147088
rect 880 146808 219120 146952
rect 880 146672 219200 146808
rect 800 145864 219200 146672
rect 880 145584 219200 145864
rect 800 145048 219200 145584
rect 800 144776 219120 145048
rect 880 144768 219120 144776
rect 880 144496 219200 144768
rect 800 143688 219200 144496
rect 880 143408 219200 143688
rect 800 143008 219200 143408
rect 800 142736 219120 143008
rect 880 142728 219120 142736
rect 880 142456 219200 142728
rect 800 141648 219200 142456
rect 880 141368 219200 141648
rect 800 140968 219200 141368
rect 800 140688 219120 140968
rect 800 140560 219200 140688
rect 880 140280 219200 140560
rect 800 139472 219200 140280
rect 880 139192 219200 139472
rect 800 138928 219200 139192
rect 800 138648 219120 138928
rect 800 138520 219200 138648
rect 880 138240 219200 138520
rect 800 137432 219200 138240
rect 880 137152 219200 137432
rect 800 136888 219200 137152
rect 800 136608 219120 136888
rect 800 136344 219200 136608
rect 880 136064 219200 136344
rect 800 135256 219200 136064
rect 880 134976 219200 135256
rect 800 134712 219200 134976
rect 800 134432 219120 134712
rect 800 134304 219200 134432
rect 880 134024 219200 134304
rect 800 133216 219200 134024
rect 880 132936 219200 133216
rect 800 132672 219200 132936
rect 800 132392 219120 132672
rect 800 132128 219200 132392
rect 880 131848 219200 132128
rect 800 131040 219200 131848
rect 880 130760 219200 131040
rect 800 130632 219200 130760
rect 800 130352 219120 130632
rect 800 130088 219200 130352
rect 880 129808 219200 130088
rect 800 129000 219200 129808
rect 880 128720 219200 129000
rect 800 128592 219200 128720
rect 800 128312 219120 128592
rect 800 127912 219200 128312
rect 880 127632 219200 127912
rect 800 126824 219200 127632
rect 880 126552 219200 126824
rect 880 126544 219120 126552
rect 800 126272 219120 126544
rect 800 125872 219200 126272
rect 880 125592 219200 125872
rect 800 124784 219200 125592
rect 880 124512 219200 124784
rect 880 124504 219120 124512
rect 800 124232 219120 124504
rect 800 123696 219200 124232
rect 880 123416 219200 123696
rect 800 122744 219200 123416
rect 880 122472 219200 122744
rect 880 122464 219120 122472
rect 800 122192 219120 122464
rect 800 121656 219200 122192
rect 880 121376 219200 121656
rect 800 120568 219200 121376
rect 880 120432 219200 120568
rect 880 120288 219120 120432
rect 800 120152 219120 120288
rect 800 119480 219200 120152
rect 880 119200 219200 119480
rect 800 118528 219200 119200
rect 880 118256 219200 118528
rect 880 118248 219120 118256
rect 800 117976 219120 118248
rect 800 117440 219200 117976
rect 880 117160 219200 117440
rect 800 116352 219200 117160
rect 880 116216 219200 116352
rect 880 116072 219120 116216
rect 800 115936 219120 116072
rect 800 115264 219200 115936
rect 880 114984 219200 115264
rect 800 114312 219200 114984
rect 880 114176 219200 114312
rect 880 114032 219120 114176
rect 800 113896 219120 114032
rect 800 113224 219200 113896
rect 880 112944 219200 113224
rect 800 112136 219200 112944
rect 880 111856 219120 112136
rect 800 111048 219200 111856
rect 880 110768 219200 111048
rect 800 110096 219200 110768
rect 880 109816 219120 110096
rect 800 109008 219200 109816
rect 880 108728 219200 109008
rect 800 108056 219200 108728
rect 800 107920 219120 108056
rect 880 107776 219120 107920
rect 880 107640 219200 107776
rect 800 106832 219200 107640
rect 880 106552 219200 106832
rect 800 106016 219200 106552
rect 800 105880 219120 106016
rect 880 105736 219120 105880
rect 880 105600 219200 105736
rect 800 104792 219200 105600
rect 880 104512 219200 104792
rect 800 103976 219200 104512
rect 800 103704 219120 103976
rect 880 103696 219120 103704
rect 880 103424 219200 103696
rect 800 102616 219200 103424
rect 880 102336 219200 102616
rect 800 101800 219200 102336
rect 800 101664 219120 101800
rect 880 101520 219120 101664
rect 880 101384 219200 101520
rect 800 100576 219200 101384
rect 880 100296 219200 100576
rect 800 99760 219200 100296
rect 800 99488 219120 99760
rect 880 99480 219120 99488
rect 880 99208 219200 99480
rect 800 98400 219200 99208
rect 880 98120 219200 98400
rect 800 97720 219200 98120
rect 800 97448 219120 97720
rect 880 97440 219120 97448
rect 880 97168 219200 97440
rect 800 96360 219200 97168
rect 880 96080 219200 96360
rect 800 95680 219200 96080
rect 800 95400 219120 95680
rect 800 95272 219200 95400
rect 880 94992 219200 95272
rect 800 94320 219200 94992
rect 880 94040 219200 94320
rect 800 93640 219200 94040
rect 800 93360 219120 93640
rect 800 93232 219200 93360
rect 880 92952 219200 93232
rect 800 92144 219200 92952
rect 880 91864 219200 92144
rect 800 91600 219200 91864
rect 800 91320 219120 91600
rect 800 91056 219200 91320
rect 880 90776 219200 91056
rect 800 90104 219200 90776
rect 880 89824 219200 90104
rect 800 89560 219200 89824
rect 800 89280 219120 89560
rect 800 89016 219200 89280
rect 880 88736 219200 89016
rect 800 87928 219200 88736
rect 880 87648 219200 87928
rect 800 87520 219200 87648
rect 800 87240 219120 87520
rect 800 86840 219200 87240
rect 880 86560 219200 86840
rect 800 85888 219200 86560
rect 880 85608 219200 85888
rect 800 85344 219200 85608
rect 800 85064 219120 85344
rect 800 84800 219200 85064
rect 880 84520 219200 84800
rect 800 83712 219200 84520
rect 880 83432 219200 83712
rect 800 83304 219200 83432
rect 800 83024 219120 83304
rect 800 82624 219200 83024
rect 880 82344 219200 82624
rect 800 81672 219200 82344
rect 880 81392 219200 81672
rect 800 81264 219200 81392
rect 800 80984 219120 81264
rect 800 80584 219200 80984
rect 880 80304 219200 80584
rect 800 79496 219200 80304
rect 880 79224 219200 79496
rect 880 79216 219120 79224
rect 800 78944 219120 79216
rect 800 78408 219200 78944
rect 880 78128 219200 78408
rect 800 77456 219200 78128
rect 880 77184 219200 77456
rect 880 77176 219120 77184
rect 800 76904 219120 77176
rect 800 76368 219200 76904
rect 880 76088 219200 76368
rect 800 75280 219200 76088
rect 880 75144 219200 75280
rect 880 75000 219120 75144
rect 800 74864 219120 75000
rect 800 74192 219200 74864
rect 880 73912 219200 74192
rect 800 73240 219200 73912
rect 880 73104 219200 73240
rect 880 72960 219120 73104
rect 800 72824 219120 72960
rect 800 72152 219200 72824
rect 880 71872 219200 72152
rect 800 71064 219200 71872
rect 880 70784 219120 71064
rect 800 69976 219200 70784
rect 880 69696 219200 69976
rect 800 69024 219200 69696
rect 880 68744 219120 69024
rect 800 67936 219200 68744
rect 880 67656 219200 67936
rect 800 66848 219200 67656
rect 880 66568 219120 66848
rect 800 65760 219200 66568
rect 880 65480 219200 65760
rect 800 64808 219200 65480
rect 880 64528 219120 64808
rect 800 63720 219200 64528
rect 880 63440 219200 63720
rect 800 62768 219200 63440
rect 800 62632 219120 62768
rect 880 62488 219120 62632
rect 880 62352 219200 62488
rect 800 61680 219200 62352
rect 880 61400 219200 61680
rect 800 60728 219200 61400
rect 800 60592 219120 60728
rect 880 60448 219120 60592
rect 880 60312 219200 60448
rect 800 59504 219200 60312
rect 880 59224 219200 59504
rect 800 58688 219200 59224
rect 800 58416 219120 58688
rect 880 58408 219120 58416
rect 880 58136 219200 58408
rect 800 57464 219200 58136
rect 880 57184 219200 57464
rect 800 56648 219200 57184
rect 800 56376 219120 56648
rect 880 56368 219120 56376
rect 880 56096 219200 56368
rect 800 55288 219200 56096
rect 880 55008 219200 55288
rect 800 54608 219200 55008
rect 800 54328 219120 54608
rect 800 54200 219200 54328
rect 880 53920 219200 54200
rect 800 53248 219200 53920
rect 880 52968 219200 53248
rect 800 52568 219200 52968
rect 800 52288 219120 52568
rect 800 52160 219200 52288
rect 880 51880 219200 52160
rect 800 51072 219200 51880
rect 880 50792 219200 51072
rect 800 50392 219200 50792
rect 800 50112 219120 50392
rect 800 49984 219200 50112
rect 880 49704 219200 49984
rect 800 49032 219200 49704
rect 880 48752 219200 49032
rect 800 48352 219200 48752
rect 800 48072 219120 48352
rect 800 47944 219200 48072
rect 880 47664 219200 47944
rect 800 46856 219200 47664
rect 880 46576 219200 46856
rect 800 46312 219200 46576
rect 800 46032 219120 46312
rect 800 45768 219200 46032
rect 880 45488 219200 45768
rect 800 44816 219200 45488
rect 880 44536 219200 44816
rect 800 44272 219200 44536
rect 800 43992 219120 44272
rect 800 43728 219200 43992
rect 880 43448 219200 43728
rect 800 42640 219200 43448
rect 880 42360 219200 42640
rect 800 42232 219200 42360
rect 800 41952 219120 42232
rect 800 41552 219200 41952
rect 880 41272 219200 41552
rect 800 40600 219200 41272
rect 880 40320 219200 40600
rect 800 40192 219200 40320
rect 800 39912 219120 40192
rect 800 39512 219200 39912
rect 880 39232 219200 39512
rect 800 38424 219200 39232
rect 880 38152 219200 38424
rect 880 38144 219120 38152
rect 800 37872 219120 38144
rect 800 37336 219200 37872
rect 880 37056 219200 37336
rect 800 36384 219200 37056
rect 880 36112 219200 36384
rect 880 36104 219120 36112
rect 800 35832 219120 36104
rect 800 35296 219200 35832
rect 880 35016 219200 35296
rect 800 34208 219200 35016
rect 880 33936 219200 34208
rect 880 33928 219120 33936
rect 800 33656 219120 33928
rect 800 33120 219200 33656
rect 880 32840 219200 33120
rect 800 32168 219200 32840
rect 880 31896 219200 32168
rect 880 31888 219120 31896
rect 800 31616 219120 31888
rect 800 31080 219200 31616
rect 880 30800 219200 31080
rect 800 29992 219200 30800
rect 880 29856 219200 29992
rect 880 29712 219120 29856
rect 800 29576 219120 29712
rect 800 29040 219200 29576
rect 880 28760 219200 29040
rect 800 27952 219200 28760
rect 880 27816 219200 27952
rect 880 27672 219120 27816
rect 800 27536 219120 27672
rect 800 26864 219200 27536
rect 880 26584 219200 26864
rect 800 25776 219200 26584
rect 880 25496 219120 25776
rect 800 24824 219200 25496
rect 880 24544 219200 24824
rect 800 23736 219200 24544
rect 880 23456 219120 23736
rect 800 22648 219200 23456
rect 880 22368 219200 22648
rect 800 21696 219200 22368
rect 800 21560 219120 21696
rect 880 21416 219120 21560
rect 880 21280 219200 21416
rect 800 20608 219200 21280
rect 880 20328 219200 20608
rect 800 19656 219200 20328
rect 800 19520 219120 19656
rect 880 19376 219120 19520
rect 880 19240 219200 19376
rect 800 18432 219200 19240
rect 880 18152 219200 18432
rect 800 17480 219200 18152
rect 800 17344 219120 17480
rect 880 17200 219120 17344
rect 880 17064 219200 17200
rect 800 16392 219200 17064
rect 880 16112 219200 16392
rect 800 15440 219200 16112
rect 800 15304 219120 15440
rect 880 15160 219120 15304
rect 880 15024 219200 15160
rect 800 14216 219200 15024
rect 880 13936 219200 14216
rect 800 13400 219200 13936
rect 800 13128 219120 13400
rect 880 13120 219120 13128
rect 880 12848 219200 13120
rect 800 12176 219200 12848
rect 880 11896 219200 12176
rect 800 11360 219200 11896
rect 800 11088 219120 11360
rect 880 11080 219120 11088
rect 880 10808 219200 11080
rect 800 10000 219200 10808
rect 880 9720 219200 10000
rect 800 9320 219200 9720
rect 800 9040 219120 9320
rect 800 8912 219200 9040
rect 880 8632 219200 8912
rect 800 7960 219200 8632
rect 880 7680 219200 7960
rect 800 7280 219200 7680
rect 800 7000 219120 7280
rect 800 6872 219200 7000
rect 880 6592 219200 6872
rect 800 5784 219200 6592
rect 880 5504 219200 5784
rect 800 5240 219200 5504
rect 800 4960 219120 5240
rect 800 4696 219200 4960
rect 880 4416 219200 4696
rect 800 3744 219200 4416
rect 880 3464 219200 3744
rect 800 3200 219200 3464
rect 800 2920 219120 3200
rect 800 2656 219200 2920
rect 880 2376 219200 2656
rect 800 1568 219200 2376
rect 880 1288 219200 1568
rect 800 1160 219200 1288
rect 800 880 219120 1160
rect 800 616 219200 880
rect 880 443 219200 616
<< metal4 >>
rect 4208 2128 4528 217648
rect 19568 2128 19888 217648
rect 34928 2128 35248 217648
rect 50288 2128 50608 217648
rect 65648 2128 65968 217648
rect 81008 2128 81328 217648
rect 96368 2128 96688 217648
rect 111728 2128 112048 217648
rect 127088 2128 127408 217648
rect 142448 2128 142768 217648
rect 157808 2128 158128 217648
rect 173168 2128 173488 217648
rect 188528 2128 188848 217648
rect 203888 2128 204208 217648
<< obsm4 >>
rect 11835 26827 19488 217157
rect 19968 26827 34848 217157
rect 35328 26827 50208 217157
rect 50688 26827 65568 217157
rect 66048 26827 80928 217157
rect 81408 26827 96288 217157
rect 96768 26827 111648 217157
rect 112128 26827 127008 217157
rect 127488 26827 142368 217157
rect 142848 26827 157728 217157
rect 158208 26827 173088 217157
rect 173568 26827 188448 217157
rect 188928 26827 203808 217157
rect 204288 26827 217797 217157
<< labels >>
rlabel metal2 s 1950 0 2006 800 6 clock
port 1 nsew signal input
rlabel metal3 s 0 3544 800 3664 6 io_dbus_addr[0]
port 2 nsew signal input
rlabel metal3 s 0 40400 800 40520 6 io_dbus_addr[10]
port 3 nsew signal input
rlabel metal3 s 0 43528 800 43648 6 io_dbus_addr[11]
port 4 nsew signal input
rlabel metal3 s 0 46656 800 46776 6 io_dbus_addr[12]
port 5 nsew signal input
rlabel metal3 s 0 49784 800 49904 6 io_dbus_addr[13]
port 6 nsew signal input
rlabel metal3 s 0 53048 800 53168 6 io_dbus_addr[14]
port 7 nsew signal input
rlabel metal3 s 0 56176 800 56296 6 io_dbus_addr[15]
port 8 nsew signal input
rlabel metal3 s 0 59304 800 59424 6 io_dbus_addr[16]
port 9 nsew signal input
rlabel metal3 s 0 62432 800 62552 6 io_dbus_addr[17]
port 10 nsew signal input
rlabel metal3 s 0 65560 800 65680 6 io_dbus_addr[18]
port 11 nsew signal input
rlabel metal3 s 0 68824 800 68944 6 io_dbus_addr[19]
port 12 nsew signal input
rlabel metal3 s 0 8712 800 8832 6 io_dbus_addr[1]
port 13 nsew signal input
rlabel metal3 s 0 71952 800 72072 6 io_dbus_addr[20]
port 14 nsew signal input
rlabel metal3 s 0 75080 800 75200 6 io_dbus_addr[21]
port 15 nsew signal input
rlabel metal3 s 0 78208 800 78328 6 io_dbus_addr[22]
port 16 nsew signal input
rlabel metal3 s 0 81472 800 81592 6 io_dbus_addr[23]
port 17 nsew signal input
rlabel metal3 s 0 84600 800 84720 6 io_dbus_addr[24]
port 18 nsew signal input
rlabel metal3 s 0 87728 800 87848 6 io_dbus_addr[25]
port 19 nsew signal input
rlabel metal3 s 0 90856 800 90976 6 io_dbus_addr[26]
port 20 nsew signal input
rlabel metal3 s 0 94120 800 94240 6 io_dbus_addr[27]
port 21 nsew signal input
rlabel metal3 s 0 97248 800 97368 6 io_dbus_addr[28]
port 22 nsew signal input
rlabel metal3 s 0 100376 800 100496 6 io_dbus_addr[29]
port 23 nsew signal input
rlabel metal3 s 0 14016 800 14136 6 io_dbus_addr[2]
port 24 nsew signal input
rlabel metal3 s 0 103504 800 103624 6 io_dbus_addr[30]
port 25 nsew signal input
rlabel metal3 s 0 106632 800 106752 6 io_dbus_addr[31]
port 26 nsew signal input
rlabel metal3 s 0 18232 800 18352 6 io_dbus_addr[3]
port 27 nsew signal input
rlabel metal3 s 0 21360 800 21480 6 io_dbus_addr[4]
port 28 nsew signal input
rlabel metal3 s 0 24624 800 24744 6 io_dbus_addr[5]
port 29 nsew signal input
rlabel metal3 s 0 27752 800 27872 6 io_dbus_addr[6]
port 30 nsew signal input
rlabel metal3 s 0 30880 800 31000 6 io_dbus_addr[7]
port 31 nsew signal input
rlabel metal3 s 0 34008 800 34128 6 io_dbus_addr[8]
port 32 nsew signal input
rlabel metal3 s 0 37136 800 37256 6 io_dbus_addr[9]
port 33 nsew signal input
rlabel metal3 s 0 4496 800 4616 6 io_dbus_ld_type[0]
port 34 nsew signal input
rlabel metal3 s 0 9800 800 9920 6 io_dbus_ld_type[1]
port 35 nsew signal input
rlabel metal3 s 0 15104 800 15224 6 io_dbus_ld_type[2]
port 36 nsew signal input
rlabel metal3 s 0 416 800 536 6 io_dbus_rd_en
port 37 nsew signal input
rlabel metal3 s 0 5584 800 5704 6 io_dbus_rdata[0]
port 38 nsew signal output
rlabel metal3 s 0 41352 800 41472 6 io_dbus_rdata[10]
port 39 nsew signal output
rlabel metal3 s 0 44616 800 44736 6 io_dbus_rdata[11]
port 40 nsew signal output
rlabel metal3 s 0 47744 800 47864 6 io_dbus_rdata[12]
port 41 nsew signal output
rlabel metal3 s 0 50872 800 50992 6 io_dbus_rdata[13]
port 42 nsew signal output
rlabel metal3 s 0 54000 800 54120 6 io_dbus_rdata[14]
port 43 nsew signal output
rlabel metal3 s 0 57264 800 57384 6 io_dbus_rdata[15]
port 44 nsew signal output
rlabel metal3 s 0 60392 800 60512 6 io_dbus_rdata[16]
port 45 nsew signal output
rlabel metal3 s 0 63520 800 63640 6 io_dbus_rdata[17]
port 46 nsew signal output
rlabel metal3 s 0 66648 800 66768 6 io_dbus_rdata[18]
port 47 nsew signal output
rlabel metal3 s 0 69776 800 69896 6 io_dbus_rdata[19]
port 48 nsew signal output
rlabel metal3 s 0 10888 800 11008 6 io_dbus_rdata[1]
port 49 nsew signal output
rlabel metal3 s 0 73040 800 73160 6 io_dbus_rdata[20]
port 50 nsew signal output
rlabel metal3 s 0 76168 800 76288 6 io_dbus_rdata[21]
port 51 nsew signal output
rlabel metal3 s 0 79296 800 79416 6 io_dbus_rdata[22]
port 52 nsew signal output
rlabel metal3 s 0 82424 800 82544 6 io_dbus_rdata[23]
port 53 nsew signal output
rlabel metal3 s 0 85688 800 85808 6 io_dbus_rdata[24]
port 54 nsew signal output
rlabel metal3 s 0 88816 800 88936 6 io_dbus_rdata[25]
port 55 nsew signal output
rlabel metal3 s 0 91944 800 92064 6 io_dbus_rdata[26]
port 56 nsew signal output
rlabel metal3 s 0 95072 800 95192 6 io_dbus_rdata[27]
port 57 nsew signal output
rlabel metal3 s 0 98200 800 98320 6 io_dbus_rdata[28]
port 58 nsew signal output
rlabel metal3 s 0 101464 800 101584 6 io_dbus_rdata[29]
port 59 nsew signal output
rlabel metal3 s 0 16192 800 16312 6 io_dbus_rdata[2]
port 60 nsew signal output
rlabel metal3 s 0 104592 800 104712 6 io_dbus_rdata[30]
port 61 nsew signal output
rlabel metal3 s 0 107720 800 107840 6 io_dbus_rdata[31]
port 62 nsew signal output
rlabel metal3 s 0 19320 800 19440 6 io_dbus_rdata[3]
port 63 nsew signal output
rlabel metal3 s 0 22448 800 22568 6 io_dbus_rdata[4]
port 64 nsew signal output
rlabel metal3 s 0 25576 800 25696 6 io_dbus_rdata[5]
port 65 nsew signal output
rlabel metal3 s 0 28840 800 28960 6 io_dbus_rdata[6]
port 66 nsew signal output
rlabel metal3 s 0 31968 800 32088 6 io_dbus_rdata[7]
port 67 nsew signal output
rlabel metal3 s 0 35096 800 35216 6 io_dbus_rdata[8]
port 68 nsew signal output
rlabel metal3 s 0 38224 800 38344 6 io_dbus_rdata[9]
port 69 nsew signal output
rlabel metal3 s 0 6672 800 6792 6 io_dbus_st_type[0]
port 70 nsew signal input
rlabel metal3 s 0 11976 800 12096 6 io_dbus_st_type[1]
port 71 nsew signal input
rlabel metal3 s 0 1368 800 1488 6 io_dbus_valid
port 72 nsew signal output
rlabel metal3 s 0 7760 800 7880 6 io_dbus_wdata[0]
port 73 nsew signal input
rlabel metal3 s 0 42440 800 42560 6 io_dbus_wdata[10]
port 74 nsew signal input
rlabel metal3 s 0 45568 800 45688 6 io_dbus_wdata[11]
port 75 nsew signal input
rlabel metal3 s 0 48832 800 48952 6 io_dbus_wdata[12]
port 76 nsew signal input
rlabel metal3 s 0 51960 800 52080 6 io_dbus_wdata[13]
port 77 nsew signal input
rlabel metal3 s 0 55088 800 55208 6 io_dbus_wdata[14]
port 78 nsew signal input
rlabel metal3 s 0 58216 800 58336 6 io_dbus_wdata[15]
port 79 nsew signal input
rlabel metal3 s 0 61480 800 61600 6 io_dbus_wdata[16]
port 80 nsew signal input
rlabel metal3 s 0 64608 800 64728 6 io_dbus_wdata[17]
port 81 nsew signal input
rlabel metal3 s 0 67736 800 67856 6 io_dbus_wdata[18]
port 82 nsew signal input
rlabel metal3 s 0 70864 800 70984 6 io_dbus_wdata[19]
port 83 nsew signal input
rlabel metal3 s 0 12928 800 13048 6 io_dbus_wdata[1]
port 84 nsew signal input
rlabel metal3 s 0 73992 800 74112 6 io_dbus_wdata[20]
port 85 nsew signal input
rlabel metal3 s 0 77256 800 77376 6 io_dbus_wdata[21]
port 86 nsew signal input
rlabel metal3 s 0 80384 800 80504 6 io_dbus_wdata[22]
port 87 nsew signal input
rlabel metal3 s 0 83512 800 83632 6 io_dbus_wdata[23]
port 88 nsew signal input
rlabel metal3 s 0 86640 800 86760 6 io_dbus_wdata[24]
port 89 nsew signal input
rlabel metal3 s 0 89904 800 90024 6 io_dbus_wdata[25]
port 90 nsew signal input
rlabel metal3 s 0 93032 800 93152 6 io_dbus_wdata[26]
port 91 nsew signal input
rlabel metal3 s 0 96160 800 96280 6 io_dbus_wdata[27]
port 92 nsew signal input
rlabel metal3 s 0 99288 800 99408 6 io_dbus_wdata[28]
port 93 nsew signal input
rlabel metal3 s 0 102416 800 102536 6 io_dbus_wdata[29]
port 94 nsew signal input
rlabel metal3 s 0 17144 800 17264 6 io_dbus_wdata[2]
port 95 nsew signal input
rlabel metal3 s 0 105680 800 105800 6 io_dbus_wdata[30]
port 96 nsew signal input
rlabel metal3 s 0 108808 800 108928 6 io_dbus_wdata[31]
port 97 nsew signal input
rlabel metal3 s 0 20408 800 20528 6 io_dbus_wdata[3]
port 98 nsew signal input
rlabel metal3 s 0 23536 800 23656 6 io_dbus_wdata[4]
port 99 nsew signal input
rlabel metal3 s 0 26664 800 26784 6 io_dbus_wdata[5]
port 100 nsew signal input
rlabel metal3 s 0 29792 800 29912 6 io_dbus_wdata[6]
port 101 nsew signal input
rlabel metal3 s 0 32920 800 33040 6 io_dbus_wdata[7]
port 102 nsew signal input
rlabel metal3 s 0 36184 800 36304 6 io_dbus_wdata[8]
port 103 nsew signal input
rlabel metal3 s 0 39312 800 39432 6 io_dbus_wdata[9]
port 104 nsew signal input
rlabel metal3 s 0 2456 800 2576 6 io_dbus_wr_en
port 105 nsew signal input
rlabel metal2 s 4250 219200 4306 220000 6 io_dmem_io_addr[0]
port 106 nsew signal output
rlabel metal2 s 11242 219200 11298 220000 6 io_dmem_io_addr[1]
port 107 nsew signal output
rlabel metal2 s 18234 219200 18290 220000 6 io_dmem_io_addr[2]
port 108 nsew signal output
rlabel metal2 s 25226 219200 25282 220000 6 io_dmem_io_addr[3]
port 109 nsew signal output
rlabel metal2 s 32218 219200 32274 220000 6 io_dmem_io_addr[4]
port 110 nsew signal output
rlabel metal2 s 37462 219200 37518 220000 6 io_dmem_io_addr[5]
port 111 nsew signal output
rlabel metal2 s 42706 219200 42762 220000 6 io_dmem_io_addr[6]
port 112 nsew signal output
rlabel metal2 s 47950 219200 48006 220000 6 io_dmem_io_addr[7]
port 113 nsew signal output
rlabel metal2 s 53194 219200 53250 220000 6 io_dmem_io_addr[8]
port 114 nsew signal output
rlabel metal2 s 846 219200 902 220000 6 io_dmem_io_cs
port 115 nsew signal output
rlabel metal2 s 5998 219200 6054 220000 6 io_dmem_io_rdata[0]
port 116 nsew signal input
rlabel metal2 s 61934 219200 61990 220000 6 io_dmem_io_rdata[10]
port 117 nsew signal input
rlabel metal2 s 65430 219200 65486 220000 6 io_dmem_io_rdata[11]
port 118 nsew signal input
rlabel metal2 s 68926 219200 68982 220000 6 io_dmem_io_rdata[12]
port 119 nsew signal input
rlabel metal2 s 72422 219200 72478 220000 6 io_dmem_io_rdata[13]
port 120 nsew signal input
rlabel metal2 s 75826 219200 75882 220000 6 io_dmem_io_rdata[14]
port 121 nsew signal input
rlabel metal2 s 79322 219200 79378 220000 6 io_dmem_io_rdata[15]
port 122 nsew signal input
rlabel metal2 s 82818 219200 82874 220000 6 io_dmem_io_rdata[16]
port 123 nsew signal input
rlabel metal2 s 86314 219200 86370 220000 6 io_dmem_io_rdata[17]
port 124 nsew signal input
rlabel metal2 s 89810 219200 89866 220000 6 io_dmem_io_rdata[18]
port 125 nsew signal input
rlabel metal2 s 93306 219200 93362 220000 6 io_dmem_io_rdata[19]
port 126 nsew signal input
rlabel metal2 s 12990 219200 13046 220000 6 io_dmem_io_rdata[1]
port 127 nsew signal input
rlabel metal2 s 96802 219200 96858 220000 6 io_dmem_io_rdata[20]
port 128 nsew signal input
rlabel metal2 s 100298 219200 100354 220000 6 io_dmem_io_rdata[21]
port 129 nsew signal input
rlabel metal2 s 103794 219200 103850 220000 6 io_dmem_io_rdata[22]
port 130 nsew signal input
rlabel metal2 s 107290 219200 107346 220000 6 io_dmem_io_rdata[23]
port 131 nsew signal input
rlabel metal2 s 110786 219200 110842 220000 6 io_dmem_io_rdata[24]
port 132 nsew signal input
rlabel metal2 s 114282 219200 114338 220000 6 io_dmem_io_rdata[25]
port 133 nsew signal input
rlabel metal2 s 117778 219200 117834 220000 6 io_dmem_io_rdata[26]
port 134 nsew signal input
rlabel metal2 s 121274 219200 121330 220000 6 io_dmem_io_rdata[27]
port 135 nsew signal input
rlabel metal2 s 124770 219200 124826 220000 6 io_dmem_io_rdata[28]
port 136 nsew signal input
rlabel metal2 s 128266 219200 128322 220000 6 io_dmem_io_rdata[29]
port 137 nsew signal input
rlabel metal2 s 19982 219200 20038 220000 6 io_dmem_io_rdata[2]
port 138 nsew signal input
rlabel metal2 s 131762 219200 131818 220000 6 io_dmem_io_rdata[30]
port 139 nsew signal input
rlabel metal2 s 135258 219200 135314 220000 6 io_dmem_io_rdata[31]
port 140 nsew signal input
rlabel metal2 s 26974 219200 27030 220000 6 io_dmem_io_rdata[3]
port 141 nsew signal input
rlabel metal2 s 33966 219200 34022 220000 6 io_dmem_io_rdata[4]
port 142 nsew signal input
rlabel metal2 s 39210 219200 39266 220000 6 io_dmem_io_rdata[5]
port 143 nsew signal input
rlabel metal2 s 44454 219200 44510 220000 6 io_dmem_io_rdata[6]
port 144 nsew signal input
rlabel metal2 s 49698 219200 49754 220000 6 io_dmem_io_rdata[7]
port 145 nsew signal input
rlabel metal2 s 54942 219200 54998 220000 6 io_dmem_io_rdata[8]
port 146 nsew signal input
rlabel metal2 s 58438 219200 58494 220000 6 io_dmem_io_rdata[9]
port 147 nsew signal input
rlabel metal2 s 7746 219200 7802 220000 6 io_dmem_io_st_type[0]
port 148 nsew signal output
rlabel metal2 s 14738 219200 14794 220000 6 io_dmem_io_st_type[1]
port 149 nsew signal output
rlabel metal2 s 21730 219200 21786 220000 6 io_dmem_io_st_type[2]
port 150 nsew signal output
rlabel metal2 s 28722 219200 28778 220000 6 io_dmem_io_st_type[3]
port 151 nsew signal output
rlabel metal2 s 9494 219200 9550 220000 6 io_dmem_io_wdata[0]
port 152 nsew signal output
rlabel metal2 s 63682 219200 63738 220000 6 io_dmem_io_wdata[10]
port 153 nsew signal output
rlabel metal2 s 67178 219200 67234 220000 6 io_dmem_io_wdata[11]
port 154 nsew signal output
rlabel metal2 s 70674 219200 70730 220000 6 io_dmem_io_wdata[12]
port 155 nsew signal output
rlabel metal2 s 74170 219200 74226 220000 6 io_dmem_io_wdata[13]
port 156 nsew signal output
rlabel metal2 s 77574 219200 77630 220000 6 io_dmem_io_wdata[14]
port 157 nsew signal output
rlabel metal2 s 81070 219200 81126 220000 6 io_dmem_io_wdata[15]
port 158 nsew signal output
rlabel metal2 s 84566 219200 84622 220000 6 io_dmem_io_wdata[16]
port 159 nsew signal output
rlabel metal2 s 88062 219200 88118 220000 6 io_dmem_io_wdata[17]
port 160 nsew signal output
rlabel metal2 s 91558 219200 91614 220000 6 io_dmem_io_wdata[18]
port 161 nsew signal output
rlabel metal2 s 95054 219200 95110 220000 6 io_dmem_io_wdata[19]
port 162 nsew signal output
rlabel metal2 s 16486 219200 16542 220000 6 io_dmem_io_wdata[1]
port 163 nsew signal output
rlabel metal2 s 98550 219200 98606 220000 6 io_dmem_io_wdata[20]
port 164 nsew signal output
rlabel metal2 s 102046 219200 102102 220000 6 io_dmem_io_wdata[21]
port 165 nsew signal output
rlabel metal2 s 105542 219200 105598 220000 6 io_dmem_io_wdata[22]
port 166 nsew signal output
rlabel metal2 s 109038 219200 109094 220000 6 io_dmem_io_wdata[23]
port 167 nsew signal output
rlabel metal2 s 112534 219200 112590 220000 6 io_dmem_io_wdata[24]
port 168 nsew signal output
rlabel metal2 s 116030 219200 116086 220000 6 io_dmem_io_wdata[25]
port 169 nsew signal output
rlabel metal2 s 119526 219200 119582 220000 6 io_dmem_io_wdata[26]
port 170 nsew signal output
rlabel metal2 s 123022 219200 123078 220000 6 io_dmem_io_wdata[27]
port 171 nsew signal output
rlabel metal2 s 126518 219200 126574 220000 6 io_dmem_io_wdata[28]
port 172 nsew signal output
rlabel metal2 s 130014 219200 130070 220000 6 io_dmem_io_wdata[29]
port 173 nsew signal output
rlabel metal2 s 23478 219200 23534 220000 6 io_dmem_io_wdata[2]
port 174 nsew signal output
rlabel metal2 s 133510 219200 133566 220000 6 io_dmem_io_wdata[30]
port 175 nsew signal output
rlabel metal2 s 137006 219200 137062 220000 6 io_dmem_io_wdata[31]
port 176 nsew signal output
rlabel metal2 s 30470 219200 30526 220000 6 io_dmem_io_wdata[3]
port 177 nsew signal output
rlabel metal2 s 35714 219200 35770 220000 6 io_dmem_io_wdata[4]
port 178 nsew signal output
rlabel metal2 s 40958 219200 41014 220000 6 io_dmem_io_wdata[5]
port 179 nsew signal output
rlabel metal2 s 46202 219200 46258 220000 6 io_dmem_io_wdata[6]
port 180 nsew signal output
rlabel metal2 s 51446 219200 51502 220000 6 io_dmem_io_wdata[7]
port 181 nsew signal output
rlabel metal2 s 56690 219200 56746 220000 6 io_dmem_io_wdata[8]
port 182 nsew signal output
rlabel metal2 s 60186 219200 60242 220000 6 io_dmem_io_wdata[9]
port 183 nsew signal output
rlabel metal2 s 2502 219200 2558 220000 6 io_dmem_io_wr_en
port 184 nsew signal output
rlabel metal3 s 0 110848 800 110968 6 io_ibus_addr[0]
port 185 nsew signal input
rlabel metal3 s 0 131928 800 132048 6 io_ibus_addr[10]
port 186 nsew signal input
rlabel metal3 s 0 134104 800 134224 6 io_ibus_addr[11]
port 187 nsew signal input
rlabel metal3 s 0 136144 800 136264 6 io_ibus_addr[12]
port 188 nsew signal input
rlabel metal3 s 0 138320 800 138440 6 io_ibus_addr[13]
port 189 nsew signal input
rlabel metal3 s 0 140360 800 140480 6 io_ibus_addr[14]
port 190 nsew signal input
rlabel metal3 s 0 142536 800 142656 6 io_ibus_addr[15]
port 191 nsew signal input
rlabel metal3 s 0 144576 800 144696 6 io_ibus_addr[16]
port 192 nsew signal input
rlabel metal3 s 0 146752 800 146872 6 io_ibus_addr[17]
port 193 nsew signal input
rlabel metal3 s 0 148792 800 148912 6 io_ibus_addr[18]
port 194 nsew signal input
rlabel metal3 s 0 150968 800 151088 6 io_ibus_addr[19]
port 195 nsew signal input
rlabel metal3 s 0 113024 800 113144 6 io_ibus_addr[1]
port 196 nsew signal input
rlabel metal3 s 0 153008 800 153128 6 io_ibus_addr[20]
port 197 nsew signal input
rlabel metal3 s 0 155184 800 155304 6 io_ibus_addr[21]
port 198 nsew signal input
rlabel metal3 s 0 157224 800 157344 6 io_ibus_addr[22]
port 199 nsew signal input
rlabel metal3 s 0 159264 800 159384 6 io_ibus_addr[23]
port 200 nsew signal input
rlabel metal3 s 0 161440 800 161560 6 io_ibus_addr[24]
port 201 nsew signal input
rlabel metal3 s 0 163480 800 163600 6 io_ibus_addr[25]
port 202 nsew signal input
rlabel metal3 s 0 165656 800 165776 6 io_ibus_addr[26]
port 203 nsew signal input
rlabel metal3 s 0 167696 800 167816 6 io_ibus_addr[27]
port 204 nsew signal input
rlabel metal3 s 0 169872 800 169992 6 io_ibus_addr[28]
port 205 nsew signal input
rlabel metal3 s 0 171912 800 172032 6 io_ibus_addr[29]
port 206 nsew signal input
rlabel metal3 s 0 115064 800 115184 6 io_ibus_addr[2]
port 207 nsew signal input
rlabel metal3 s 0 174088 800 174208 6 io_ibus_addr[30]
port 208 nsew signal input
rlabel metal3 s 0 176128 800 176248 6 io_ibus_addr[31]
port 209 nsew signal input
rlabel metal3 s 0 117240 800 117360 6 io_ibus_addr[3]
port 210 nsew signal input
rlabel metal3 s 0 119280 800 119400 6 io_ibus_addr[4]
port 211 nsew signal input
rlabel metal3 s 0 121456 800 121576 6 io_ibus_addr[5]
port 212 nsew signal input
rlabel metal3 s 0 123496 800 123616 6 io_ibus_addr[6]
port 213 nsew signal input
rlabel metal3 s 0 125672 800 125792 6 io_ibus_addr[7]
port 214 nsew signal input
rlabel metal3 s 0 127712 800 127832 6 io_ibus_addr[8]
port 215 nsew signal input
rlabel metal3 s 0 129888 800 130008 6 io_ibus_addr[9]
port 216 nsew signal input
rlabel metal3 s 0 111936 800 112056 6 io_ibus_inst[0]
port 217 nsew signal output
rlabel metal3 s 0 133016 800 133136 6 io_ibus_inst[10]
port 218 nsew signal output
rlabel metal3 s 0 135056 800 135176 6 io_ibus_inst[11]
port 219 nsew signal output
rlabel metal3 s 0 137232 800 137352 6 io_ibus_inst[12]
port 220 nsew signal output
rlabel metal3 s 0 139272 800 139392 6 io_ibus_inst[13]
port 221 nsew signal output
rlabel metal3 s 0 141448 800 141568 6 io_ibus_inst[14]
port 222 nsew signal output
rlabel metal3 s 0 143488 800 143608 6 io_ibus_inst[15]
port 223 nsew signal output
rlabel metal3 s 0 145664 800 145784 6 io_ibus_inst[16]
port 224 nsew signal output
rlabel metal3 s 0 147704 800 147824 6 io_ibus_inst[17]
port 225 nsew signal output
rlabel metal3 s 0 149880 800 150000 6 io_ibus_inst[18]
port 226 nsew signal output
rlabel metal3 s 0 151920 800 152040 6 io_ibus_inst[19]
port 227 nsew signal output
rlabel metal3 s 0 114112 800 114232 6 io_ibus_inst[1]
port 228 nsew signal output
rlabel metal3 s 0 154096 800 154216 6 io_ibus_inst[20]
port 229 nsew signal output
rlabel metal3 s 0 156136 800 156256 6 io_ibus_inst[21]
port 230 nsew signal output
rlabel metal3 s 0 158312 800 158432 6 io_ibus_inst[22]
port 231 nsew signal output
rlabel metal3 s 0 160352 800 160472 6 io_ibus_inst[23]
port 232 nsew signal output
rlabel metal3 s 0 162528 800 162648 6 io_ibus_inst[24]
port 233 nsew signal output
rlabel metal3 s 0 164568 800 164688 6 io_ibus_inst[25]
port 234 nsew signal output
rlabel metal3 s 0 166744 800 166864 6 io_ibus_inst[26]
port 235 nsew signal output
rlabel metal3 s 0 168784 800 168904 6 io_ibus_inst[27]
port 236 nsew signal output
rlabel metal3 s 0 170960 800 171080 6 io_ibus_inst[28]
port 237 nsew signal output
rlabel metal3 s 0 173000 800 173120 6 io_ibus_inst[29]
port 238 nsew signal output
rlabel metal3 s 0 116152 800 116272 6 io_ibus_inst[2]
port 239 nsew signal output
rlabel metal3 s 0 175176 800 175296 6 io_ibus_inst[30]
port 240 nsew signal output
rlabel metal3 s 0 177216 800 177336 6 io_ibus_inst[31]
port 241 nsew signal output
rlabel metal3 s 0 118328 800 118448 6 io_ibus_inst[3]
port 242 nsew signal output
rlabel metal3 s 0 120368 800 120488 6 io_ibus_inst[4]
port 243 nsew signal output
rlabel metal3 s 0 122544 800 122664 6 io_ibus_inst[5]
port 244 nsew signal output
rlabel metal3 s 0 124584 800 124704 6 io_ibus_inst[6]
port 245 nsew signal output
rlabel metal3 s 0 126624 800 126744 6 io_ibus_inst[7]
port 246 nsew signal output
rlabel metal3 s 0 128800 800 128920 6 io_ibus_inst[8]
port 247 nsew signal output
rlabel metal3 s 0 130840 800 130960 6 io_ibus_inst[9]
port 248 nsew signal output
rlabel metal3 s 0 109896 800 110016 6 io_ibus_valid
port 249 nsew signal output
rlabel metal2 s 29918 0 29974 800 6 io_imem_io_addr[0]
port 250 nsew signal output
rlabel metal3 s 219200 132472 220000 132592 6 io_imem_io_addr[1]
port 251 nsew signal output
rlabel metal2 s 149150 219200 149206 220000 6 io_imem_io_addr[2]
port 252 nsew signal output
rlabel metal2 s 150898 219200 150954 220000 6 io_imem_io_addr[3]
port 253 nsew signal output
rlabel metal2 s 53930 0 53986 800 6 io_imem_io_addr[4]
port 254 nsew signal output
rlabel metal2 s 65890 0 65946 800 6 io_imem_io_addr[5]
port 255 nsew signal output
rlabel metal2 s 77850 0 77906 800 6 io_imem_io_addr[6]
port 256 nsew signal output
rlabel metal2 s 89902 0 89958 800 6 io_imem_io_addr[7]
port 257 nsew signal output
rlabel metal3 s 219200 155184 220000 155304 6 io_imem_io_addr[8]
port 258 nsew signal output
rlabel metal3 s 219200 120232 220000 120352 6 io_imem_io_cs
port 259 nsew signal output
rlabel metal2 s 140502 219200 140558 220000 6 io_imem_io_rdata[0]
port 260 nsew signal input
rlabel metal3 s 219200 163344 220000 163464 6 io_imem_io_rdata[10]
port 261 nsew signal input
rlabel metal3 s 0 192992 800 193112 6 io_imem_io_rdata[11]
port 262 nsew signal input
rlabel metal3 s 219200 169464 220000 169584 6 io_imem_io_rdata[12]
port 263 nsew signal input
rlabel metal3 s 219200 173680 220000 173800 6 io_imem_io_rdata[13]
port 264 nsew signal input
rlabel metal2 s 121918 0 121974 800 6 io_imem_io_rdata[14]
port 265 nsew signal input
rlabel metal2 s 129922 0 129978 800 6 io_imem_io_rdata[15]
port 266 nsew signal input
rlabel metal2 s 137926 0 137982 800 6 io_imem_io_rdata[16]
port 267 nsew signal input
rlabel metal3 s 0 201424 800 201544 6 io_imem_io_rdata[17]
port 268 nsew signal input
rlabel metal3 s 0 203600 800 203720 6 io_imem_io_rdata[18]
port 269 nsew signal input
rlabel metal2 s 192850 219200 192906 220000 6 io_imem_io_rdata[19]
port 270 nsew signal input
rlabel metal2 s 145746 219200 145802 220000 6 io_imem_io_rdata[1]
port 271 nsew signal input
rlabel metal3 s 0 206728 800 206848 6 io_imem_io_rdata[20]
port 272 nsew signal input
rlabel metal2 s 165894 0 165950 800 6 io_imem_io_rdata[21]
port 273 nsew signal input
rlabel metal2 s 199842 219200 199898 220000 6 io_imem_io_rdata[22]
port 274 nsew signal input
rlabel metal3 s 0 209856 800 209976 6 io_imem_io_rdata[23]
port 275 nsew signal input
rlabel metal3 s 0 212032 800 212152 6 io_imem_io_rdata[24]
port 276 nsew signal input
rlabel metal3 s 219200 198296 220000 198416 6 io_imem_io_rdata[25]
port 277 nsew signal input
rlabel metal2 s 205086 219200 205142 220000 6 io_imem_io_rdata[26]
port 278 nsew signal input
rlabel metal2 s 206834 219200 206890 220000 6 io_imem_io_rdata[27]
port 279 nsew signal input
rlabel metal2 s 193862 0 193918 800 6 io_imem_io_rdata[28]
port 280 nsew signal input
rlabel metal2 s 213826 219200 213882 220000 6 io_imem_io_rdata[29]
port 281 nsew signal input
rlabel metal2 s 37922 0 37978 800 6 io_imem_io_rdata[2]
port 282 nsew signal input
rlabel metal3 s 219200 212712 220000 212832 6 io_imem_io_rdata[30]
port 283 nsew signal input
rlabel metal3 s 219200 214752 220000 214872 6 io_imem_io_rdata[31]
port 284 nsew signal input
rlabel metal2 s 49882 0 49938 800 6 io_imem_io_rdata[3]
port 285 nsew signal input
rlabel metal3 s 0 187824 800 187944 6 io_imem_io_rdata[4]
port 286 nsew signal input
rlabel metal3 s 0 188776 800 188896 6 io_imem_io_rdata[5]
port 287 nsew signal input
rlabel metal3 s 219200 146888 220000 147008 6 io_imem_io_rdata[6]
port 288 nsew signal input
rlabel metal3 s 219200 150968 220000 151088 6 io_imem_io_rdata[7]
port 289 nsew signal input
rlabel metal2 s 168378 219200 168434 220000 6 io_imem_io_rdata[8]
port 290 nsew signal input
rlabel metal3 s 0 190952 800 191072 6 io_imem_io_rdata[9]
port 291 nsew signal input
rlabel metal3 s 219200 128392 220000 128512 6 io_imem_io_st_type[0]
port 292 nsew signal output
rlabel metal2 s 147494 219200 147550 220000 6 io_imem_io_st_type[1]
port 293 nsew signal output
rlabel metal2 s 41878 0 41934 800 6 io_imem_io_st_type[2]
port 294 nsew signal output
rlabel metal2 s 152646 219200 152702 220000 6 io_imem_io_st_type[3]
port 295 nsew signal output
rlabel metal2 s 142250 219200 142306 220000 6 io_imem_io_wdata[0]
port 296 nsew signal output
rlabel metal3 s 219200 165384 220000 165504 6 io_imem_io_wdata[10]
port 297 nsew signal output
rlabel metal2 s 113914 0 113970 800 6 io_imem_io_wdata[11]
port 298 nsew signal output
rlabel metal3 s 0 195168 800 195288 6 io_imem_io_wdata[12]
port 299 nsew signal output
rlabel metal3 s 219200 175720 220000 175840 6 io_imem_io_wdata[13]
port 300 nsew signal output
rlabel metal2 s 125874 0 125930 800 6 io_imem_io_wdata[14]
port 301 nsew signal output
rlabel metal2 s 133878 0 133934 800 6 io_imem_io_wdata[15]
port 302 nsew signal output
rlabel metal2 s 141882 0 141938 800 6 io_imem_io_wdata[16]
port 303 nsew signal output
rlabel metal2 s 189354 219200 189410 220000 6 io_imem_io_wdata[17]
port 304 nsew signal output
rlabel metal2 s 149886 0 149942 800 6 io_imem_io_wdata[18]
port 305 nsew signal output
rlabel metal2 s 194598 219200 194654 220000 6 io_imem_io_wdata[19]
port 306 nsew signal output
rlabel metal3 s 0 185648 800 185768 6 io_imem_io_wdata[1]
port 307 nsew signal output
rlabel metal2 s 161846 0 161902 800 6 io_imem_io_wdata[20]
port 308 nsew signal output
rlabel metal3 s 219200 185920 220000 186040 6 io_imem_io_wdata[21]
port 309 nsew signal output
rlabel metal3 s 219200 188096 220000 188216 6 io_imem_io_wdata[22]
port 310 nsew signal output
rlabel metal3 s 219200 194216 220000 194336 6 io_imem_io_wdata[23]
port 311 nsew signal output
rlabel metal3 s 219200 196256 220000 196376 6 io_imem_io_wdata[24]
port 312 nsew signal output
rlabel metal3 s 219200 200336 220000 200456 6 io_imem_io_wdata[25]
port 313 nsew signal output
rlabel metal2 s 185858 0 185914 800 6 io_imem_io_wdata[26]
port 314 nsew signal output
rlabel metal2 s 189906 0 189962 800 6 io_imem_io_wdata[27]
port 315 nsew signal output
rlabel metal2 s 197910 0 197966 800 6 io_imem_io_wdata[28]
port 316 nsew signal output
rlabel metal3 s 0 218288 800 218408 6 io_imem_io_wdata[29]
port 317 nsew signal output
rlabel metal2 s 45926 0 45982 800 6 io_imem_io_wdata[2]
port 318 nsew signal output
rlabel metal2 s 219070 219200 219126 220000 6 io_imem_io_wdata[30]
port 319 nsew signal output
rlabel metal2 s 213918 0 213974 800 6 io_imem_io_wdata[31]
port 320 nsew signal output
rlabel metal2 s 154394 219200 154450 220000 6 io_imem_io_wdata[3]
port 321 nsew signal output
rlabel metal2 s 57886 0 57942 800 6 io_imem_io_wdata[4]
port 322 nsew signal output
rlabel metal2 s 69938 0 69994 800 6 io_imem_io_wdata[5]
port 323 nsew signal output
rlabel metal2 s 81898 0 81954 800 6 io_imem_io_wdata[6]
port 324 nsew signal output
rlabel metal2 s 166630 219200 166686 220000 6 io_imem_io_wdata[7]
port 325 nsew signal output
rlabel metal3 s 219200 157224 220000 157344 6 io_imem_io_wdata[8]
port 326 nsew signal output
rlabel metal2 s 170126 219200 170182 220000 6 io_imem_io_wdata[9]
port 327 nsew signal output
rlabel metal3 s 219200 122272 220000 122392 6 io_imem_io_wr_en
port 328 nsew signal output
rlabel metal3 s 219200 124312 220000 124432 6 io_m1_ack_i
port 329 nsew signal input
rlabel metal2 s 17866 0 17922 800 6 io_m1_addr_sel
port 330 nsew signal output
rlabel metal3 s 0 184560 800 184680 6 io_m1_data_i[0]
port 331 nsew signal input
rlabel metal2 s 105910 0 105966 800 6 io_m1_data_i[10]
port 332 nsew signal input
rlabel metal3 s 0 194080 800 194200 6 io_m1_data_i[11]
port 333 nsew signal input
rlabel metal2 s 177118 219200 177174 220000 6 io_m1_data_i[12]
port 334 nsew signal input
rlabel metal3 s 0 196120 800 196240 6 io_m1_data_i[13]
port 335 nsew signal input
rlabel metal2 s 182362 219200 182418 220000 6 io_m1_data_i[14]
port 336 nsew signal input
rlabel metal3 s 0 198296 800 198416 6 io_m1_data_i[15]
port 337 nsew signal input
rlabel metal2 s 187606 219200 187662 220000 6 io_m1_data_i[16]
port 338 nsew signal input
rlabel metal3 s 0 202512 800 202632 6 io_m1_data_i[17]
port 339 nsew signal input
rlabel metal2 s 153842 0 153898 800 6 io_m1_data_i[18]
port 340 nsew signal input
rlabel metal2 s 196346 219200 196402 220000 6 io_m1_data_i[19]
port 341 nsew signal input
rlabel metal2 s 33874 0 33930 800 6 io_m1_data_i[1]
port 342 nsew signal input
rlabel metal3 s 0 207816 800 207936 6 io_m1_data_i[20]
port 343 nsew signal input
rlabel metal2 s 169850 0 169906 800 6 io_m1_data_i[21]
port 344 nsew signal input
rlabel metal3 s 219200 190136 220000 190256 6 io_m1_data_i[22]
port 345 nsew signal input
rlabel metal2 s 173898 0 173954 800 6 io_m1_data_i[23]
port 346 nsew signal input
rlabel metal2 s 177854 0 177910 800 6 io_m1_data_i[24]
port 347 nsew signal input
rlabel metal3 s 0 214072 800 214192 6 io_m1_data_i[25]
port 348 nsew signal input
rlabel metal3 s 0 217200 800 217320 6 io_m1_data_i[26]
port 349 nsew signal input
rlabel metal2 s 208582 219200 208638 220000 6 io_m1_data_i[27]
port 350 nsew signal input
rlabel metal2 s 212078 219200 212134 220000 6 io_m1_data_i[28]
port 351 nsew signal input
rlabel metal2 s 215574 219200 215630 220000 6 io_m1_data_i[29]
port 352 nsew signal input
rlabel metal3 s 219200 136688 220000 136808 6 io_m1_data_i[2]
port 353 nsew signal input
rlabel metal3 s 0 219376 800 219496 6 io_m1_data_i[30]
port 354 nsew signal input
rlabel metal3 s 219200 216792 220000 216912 6 io_m1_data_i[31]
port 355 nsew signal input
rlabel metal2 s 156142 219200 156198 220000 6 io_m1_data_i[3]
port 356 nsew signal input
rlabel metal3 s 219200 142808 220000 142928 6 io_m1_data_i[4]
port 357 nsew signal input
rlabel metal2 s 161386 219200 161442 220000 6 io_m1_data_i[5]
port 358 nsew signal input
rlabel metal2 s 164882 219200 164938 220000 6 io_m1_data_i[6]
port 359 nsew signal input
rlabel metal3 s 219200 153008 220000 153128 6 io_m1_data_i[7]
port 360 nsew signal input
rlabel metal3 s 0 189864 800 189984 6 io_m1_data_i[8]
port 361 nsew signal input
rlabel metal3 s 0 191904 800 192024 6 io_m1_data_i[9]
port 362 nsew signal input
rlabel metal2 s 21914 0 21970 800 6 io_m2_ack_i
port 363 nsew signal input
rlabel metal2 s 25870 0 25926 800 6 io_m2_addr_sel
port 364 nsew signal output
rlabel metal2 s 143998 219200 144054 220000 6 io_m2_data_i[0]
port 365 nsew signal input
rlabel metal2 s 109866 0 109922 800 6 io_m2_data_i[10]
port 366 nsew signal input
rlabel metal2 s 173622 219200 173678 220000 6 io_m2_data_i[11]
port 367 nsew signal input
rlabel metal2 s 178866 219200 178922 220000 6 io_m2_data_i[12]
port 368 nsew signal input
rlabel metal2 s 180614 219200 180670 220000 6 io_m2_data_i[13]
port 369 nsew signal input
rlabel metal3 s 0 197208 800 197328 6 io_m2_data_i[14]
port 370 nsew signal input
rlabel metal3 s 0 199384 800 199504 6 io_m2_data_i[15]
port 371 nsew signal input
rlabel metal2 s 145930 0 145986 800 6 io_m2_data_i[16]
port 372 nsew signal input
rlabel metal3 s 219200 177760 220000 177880 6 io_m2_data_i[17]
port 373 nsew signal input
rlabel metal2 s 191102 219200 191158 220000 6 io_m2_data_i[18]
port 374 nsew signal input
rlabel metal3 s 0 204552 800 204672 6 io_m2_data_i[19]
port 375 nsew signal input
rlabel metal3 s 219200 134512 220000 134632 6 io_m2_data_i[1]
port 376 nsew signal input
rlabel metal3 s 219200 181840 220000 181960 6 io_m2_data_i[20]
port 377 nsew signal input
rlabel metal3 s 0 208768 800 208888 6 io_m2_data_i[21]
port 378 nsew signal input
rlabel metal2 s 201590 219200 201646 220000 6 io_m2_data_i[22]
port 379 nsew signal input
rlabel metal3 s 0 210944 800 211064 6 io_m2_data_i[23]
port 380 nsew signal input
rlabel metal2 s 181902 0 181958 800 6 io_m2_data_i[24]
port 381 nsew signal input
rlabel metal3 s 0 215160 800 215280 6 io_m2_data_i[25]
port 382 nsew signal input
rlabel metal3 s 219200 202376 220000 202496 6 io_m2_data_i[26]
port 383 nsew signal input
rlabel metal3 s 219200 206592 220000 206712 6 io_m2_data_i[27]
port 384 nsew signal input
rlabel metal3 s 219200 208632 220000 208752 6 io_m2_data_i[28]
port 385 nsew signal input
rlabel metal2 s 201866 0 201922 800 6 io_m2_data_i[29]
port 386 nsew signal input
rlabel metal3 s 219200 138728 220000 138848 6 io_m2_data_i[2]
port 387 nsew signal input
rlabel metal2 s 205914 0 205970 800 6 io_m2_data_i[30]
port 388 nsew signal input
rlabel metal2 s 217874 0 217930 800 6 io_m2_data_i[31]
port 389 nsew signal input
rlabel metal2 s 157890 219200 157946 220000 6 io_m2_data_i[3]
port 390 nsew signal input
rlabel metal3 s 219200 144848 220000 144968 6 io_m2_data_i[4]
port 391 nsew signal input
rlabel metal2 s 73894 0 73950 800 6 io_m2_data_i[5]
port 392 nsew signal input
rlabel metal3 s 219200 148928 220000 149048 6 io_m2_data_i[6]
port 393 nsew signal input
rlabel metal2 s 93858 0 93914 800 6 io_m2_data_i[7]
port 394 nsew signal input
rlabel metal3 s 219200 159264 220000 159384 6 io_m2_data_i[8]
port 395 nsew signal input
rlabel metal3 s 219200 161304 220000 161424 6 io_m2_data_i[9]
port 396 nsew signal input
rlabel metal3 s 0 180344 800 180464 6 io_m3_ack_i
port 397 nsew signal input
rlabel metal3 s 0 181432 800 181552 6 io_m3_addr_sel
port 398 nsew signal output
rlabel metal3 s 219200 130432 220000 130552 6 io_m3_data_i[0]
port 399 nsew signal input
rlabel metal3 s 219200 167424 220000 167544 6 io_m3_data_i[10]
port 400 nsew signal input
rlabel metal2 s 175370 219200 175426 220000 6 io_m3_data_i[11]
port 401 nsew signal input
rlabel metal3 s 219200 171640 220000 171760 6 io_m3_data_i[12]
port 402 nsew signal input
rlabel metal2 s 117870 0 117926 800 6 io_m3_data_i[13]
port 403 nsew signal input
rlabel metal2 s 184110 219200 184166 220000 6 io_m3_data_i[14]
port 404 nsew signal input
rlabel metal2 s 185858 219200 185914 220000 6 io_m3_data_i[15]
port 405 nsew signal input
rlabel metal3 s 0 200336 800 200456 6 io_m3_data_i[16]
port 406 nsew signal input
rlabel metal3 s 219200 179800 220000 179920 6 io_m3_data_i[17]
port 407 nsew signal input
rlabel metal2 s 157890 0 157946 800 6 io_m3_data_i[18]
port 408 nsew signal input
rlabel metal3 s 0 205640 800 205760 6 io_m3_data_i[19]
port 409 nsew signal input
rlabel metal3 s 0 186736 800 186856 6 io_m3_data_i[1]
port 410 nsew signal input
rlabel metal3 s 219200 183880 220000 184000 6 io_m3_data_i[20]
port 411 nsew signal input
rlabel metal2 s 198094 219200 198150 220000 6 io_m3_data_i[21]
port 412 nsew signal input
rlabel metal3 s 219200 192176 220000 192296 6 io_m3_data_i[22]
port 413 nsew signal input
rlabel metal2 s 203338 219200 203394 220000 6 io_m3_data_i[23]
port 414 nsew signal input
rlabel metal3 s 0 212984 800 213104 6 io_m3_data_i[24]
port 415 nsew signal input
rlabel metal3 s 0 216248 800 216368 6 io_m3_data_i[25]
port 416 nsew signal input
rlabel metal3 s 219200 204552 220000 204672 6 io_m3_data_i[26]
port 417 nsew signal input
rlabel metal2 s 210330 219200 210386 220000 6 io_m3_data_i[27]
port 418 nsew signal input
rlabel metal3 s 219200 210672 220000 210792 6 io_m3_data_i[28]
port 419 nsew signal input
rlabel metal2 s 217322 219200 217378 220000 6 io_m3_data_i[29]
port 420 nsew signal input
rlabel metal3 s 219200 140768 220000 140888 6 io_m3_data_i[2]
port 421 nsew signal input
rlabel metal2 s 209870 0 209926 800 6 io_m3_data_i[30]
port 422 nsew signal input
rlabel metal3 s 219200 218832 220000 218952 6 io_m3_data_i[31]
port 423 nsew signal input
rlabel metal2 s 159638 219200 159694 220000 6 io_m3_data_i[3]
port 424 nsew signal input
rlabel metal2 s 61934 0 61990 800 6 io_m3_data_i[4]
port 425 nsew signal input
rlabel metal2 s 163134 219200 163190 220000 6 io_m3_data_i[5]
port 426 nsew signal input
rlabel metal2 s 85854 0 85910 800 6 io_m3_data_i[6]
port 427 nsew signal input
rlabel metal2 s 97906 0 97962 800 6 io_m3_data_i[7]
port 428 nsew signal input
rlabel metal2 s 101862 0 101918 800 6 io_m3_data_i[8]
port 429 nsew signal input
rlabel metal2 s 171874 219200 171930 220000 6 io_m3_data_i[9]
port 430 nsew signal input
rlabel metal3 s 219200 111936 220000 112056 6 io_spi_clk
port 431 nsew signal output
rlabel metal2 s 138754 219200 138810 220000 6 io_spi_clk_en
port 432 nsew signal output
rlabel metal3 s 219200 113976 220000 114096 6 io_spi_cs
port 433 nsew signal output
rlabel metal3 s 0 182520 800 182640 6 io_spi_cs_en
port 434 nsew signal output
rlabel metal3 s 0 178304 800 178424 6 io_spi_irq
port 435 nsew signal output
rlabel metal2 s 9862 0 9918 800 6 io_spi_miso
port 436 nsew signal input
rlabel metal3 s 219200 116016 220000 116136 6 io_spi_mosi
port 437 nsew signal output
rlabel metal3 s 219200 126352 220000 126472 6 io_spi_mosi_en
port 438 nsew signal output
rlabel metal3 s 0 179392 800 179512 6 io_uart_irq
port 439 nsew signal output
rlabel metal2 s 13910 0 13966 800 6 io_uart_rx
port 440 nsew signal input
rlabel metal3 s 219200 118056 220000 118176 6 io_uart_tx
port 441 nsew signal output
rlabel metal3 s 0 183608 800 183728 6 io_uart_tx_en
port 442 nsew signal output
rlabel metal3 s 219200 5040 220000 5160 6 io_wbm_m2s_addr[0]
port 443 nsew signal output
rlabel metal3 s 219200 54408 220000 54528 6 io_wbm_m2s_addr[10]
port 444 nsew signal output
rlabel metal3 s 219200 58488 220000 58608 6 io_wbm_m2s_addr[11]
port 445 nsew signal output
rlabel metal3 s 219200 62568 220000 62688 6 io_wbm_m2s_addr[12]
port 446 nsew signal output
rlabel metal3 s 219200 66648 220000 66768 6 io_wbm_m2s_addr[13]
port 447 nsew signal output
rlabel metal3 s 219200 70864 220000 70984 6 io_wbm_m2s_addr[14]
port 448 nsew signal output
rlabel metal3 s 219200 74944 220000 75064 6 io_wbm_m2s_addr[15]
port 449 nsew signal output
rlabel metal3 s 219200 11160 220000 11280 6 io_wbm_m2s_addr[1]
port 450 nsew signal output
rlabel metal3 s 219200 17280 220000 17400 6 io_wbm_m2s_addr[2]
port 451 nsew signal output
rlabel metal3 s 219200 23536 220000 23656 6 io_wbm_m2s_addr[3]
port 452 nsew signal output
rlabel metal3 s 219200 29656 220000 29776 6 io_wbm_m2s_addr[4]
port 453 nsew signal output
rlabel metal3 s 219200 33736 220000 33856 6 io_wbm_m2s_addr[5]
port 454 nsew signal output
rlabel metal3 s 219200 37952 220000 38072 6 io_wbm_m2s_addr[6]
port 455 nsew signal output
rlabel metal3 s 219200 42032 220000 42152 6 io_wbm_m2s_addr[7]
port 456 nsew signal output
rlabel metal3 s 219200 46112 220000 46232 6 io_wbm_m2s_addr[8]
port 457 nsew signal output
rlabel metal3 s 219200 50192 220000 50312 6 io_wbm_m2s_addr[9]
port 458 nsew signal output
rlabel metal3 s 219200 7080 220000 7200 6 io_wbm_m2s_data[0]
port 459 nsew signal output
rlabel metal3 s 219200 56448 220000 56568 6 io_wbm_m2s_data[10]
port 460 nsew signal output
rlabel metal3 s 219200 60528 220000 60648 6 io_wbm_m2s_data[11]
port 461 nsew signal output
rlabel metal3 s 219200 64608 220000 64728 6 io_wbm_m2s_data[12]
port 462 nsew signal output
rlabel metal3 s 219200 68824 220000 68944 6 io_wbm_m2s_data[13]
port 463 nsew signal output
rlabel metal3 s 219200 72904 220000 73024 6 io_wbm_m2s_data[14]
port 464 nsew signal output
rlabel metal3 s 219200 76984 220000 77104 6 io_wbm_m2s_data[15]
port 465 nsew signal output
rlabel metal3 s 219200 79024 220000 79144 6 io_wbm_m2s_data[16]
port 466 nsew signal output
rlabel metal3 s 219200 81064 220000 81184 6 io_wbm_m2s_data[17]
port 467 nsew signal output
rlabel metal3 s 219200 83104 220000 83224 6 io_wbm_m2s_data[18]
port 468 nsew signal output
rlabel metal3 s 219200 85144 220000 85264 6 io_wbm_m2s_data[19]
port 469 nsew signal output
rlabel metal3 s 219200 13200 220000 13320 6 io_wbm_m2s_data[1]
port 470 nsew signal output
rlabel metal3 s 219200 87320 220000 87440 6 io_wbm_m2s_data[20]
port 471 nsew signal output
rlabel metal3 s 219200 89360 220000 89480 6 io_wbm_m2s_data[21]
port 472 nsew signal output
rlabel metal3 s 219200 91400 220000 91520 6 io_wbm_m2s_data[22]
port 473 nsew signal output
rlabel metal3 s 219200 93440 220000 93560 6 io_wbm_m2s_data[23]
port 474 nsew signal output
rlabel metal3 s 219200 95480 220000 95600 6 io_wbm_m2s_data[24]
port 475 nsew signal output
rlabel metal3 s 219200 97520 220000 97640 6 io_wbm_m2s_data[25]
port 476 nsew signal output
rlabel metal3 s 219200 99560 220000 99680 6 io_wbm_m2s_data[26]
port 477 nsew signal output
rlabel metal3 s 219200 101600 220000 101720 6 io_wbm_m2s_data[27]
port 478 nsew signal output
rlabel metal3 s 219200 103776 220000 103896 6 io_wbm_m2s_data[28]
port 479 nsew signal output
rlabel metal3 s 219200 105816 220000 105936 6 io_wbm_m2s_data[29]
port 480 nsew signal output
rlabel metal3 s 219200 19456 220000 19576 6 io_wbm_m2s_data[2]
port 481 nsew signal output
rlabel metal3 s 219200 107856 220000 107976 6 io_wbm_m2s_data[30]
port 482 nsew signal output
rlabel metal3 s 219200 109896 220000 110016 6 io_wbm_m2s_data[31]
port 483 nsew signal output
rlabel metal3 s 219200 25576 220000 25696 6 io_wbm_m2s_data[3]
port 484 nsew signal output
rlabel metal3 s 219200 31696 220000 31816 6 io_wbm_m2s_data[4]
port 485 nsew signal output
rlabel metal3 s 219200 35912 220000 36032 6 io_wbm_m2s_data[5]
port 486 nsew signal output
rlabel metal3 s 219200 39992 220000 40112 6 io_wbm_m2s_data[6]
port 487 nsew signal output
rlabel metal3 s 219200 44072 220000 44192 6 io_wbm_m2s_data[7]
port 488 nsew signal output
rlabel metal3 s 219200 48152 220000 48272 6 io_wbm_m2s_data[8]
port 489 nsew signal output
rlabel metal3 s 219200 52368 220000 52488 6 io_wbm_m2s_data[9]
port 490 nsew signal output
rlabel metal3 s 219200 9120 220000 9240 6 io_wbm_m2s_sel[0]
port 491 nsew signal output
rlabel metal3 s 219200 15240 220000 15360 6 io_wbm_m2s_sel[1]
port 492 nsew signal output
rlabel metal3 s 219200 21496 220000 21616 6 io_wbm_m2s_sel[2]
port 493 nsew signal output
rlabel metal3 s 219200 27616 220000 27736 6 io_wbm_m2s_sel[3]
port 494 nsew signal output
rlabel metal3 s 219200 960 220000 1080 6 io_wbm_m2s_stb
port 495 nsew signal output
rlabel metal3 s 219200 3000 220000 3120 6 io_wbm_m2s_we
port 496 nsew signal output
rlabel metal2 s 5906 0 5962 800 6 reset
port 497 nsew signal input
rlabel metal4 s 4208 2128 4528 217648 6 vccd1
port 498 nsew power input
rlabel metal4 s 34928 2128 35248 217648 6 vccd1
port 498 nsew power input
rlabel metal4 s 65648 2128 65968 217648 6 vccd1
port 498 nsew power input
rlabel metal4 s 96368 2128 96688 217648 6 vccd1
port 498 nsew power input
rlabel metal4 s 127088 2128 127408 217648 6 vccd1
port 498 nsew power input
rlabel metal4 s 157808 2128 158128 217648 6 vccd1
port 498 nsew power input
rlabel metal4 s 188528 2128 188848 217648 6 vccd1
port 498 nsew power input
rlabel metal4 s 19568 2128 19888 217648 6 vssd1
port 499 nsew ground input
rlabel metal4 s 50288 2128 50608 217648 6 vssd1
port 499 nsew ground input
rlabel metal4 s 81008 2128 81328 217648 6 vssd1
port 499 nsew ground input
rlabel metal4 s 111728 2128 112048 217648 6 vssd1
port 499 nsew ground input
rlabel metal4 s 142448 2128 142768 217648 6 vssd1
port 499 nsew ground input
rlabel metal4 s 173168 2128 173488 217648 6 vssd1
port 499 nsew ground input
rlabel metal4 s 203888 2128 204208 217648 6 vssd1
port 499 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 220000 220000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 19420490
string GDS_FILE /home/ali112000/Desktop/mpw/UETRV-ECORE/openlane/Wishbone_InterConnect/runs/Wishbone_InterConnect/results/finishing/WB_InterConnect.magic.gds
string GDS_START 1020738
<< end >>

