magic
tech sky130A
magscale 1 2
timestamp 1647675757
<< obsli1 >>
rect 1104 2159 78844 77809
<< obsm1 >>
rect 1104 2128 78844 77920
<< metal2 >>
rect 1398 79200 1454 80000
rect 4158 79200 4214 80000
rect 6918 79200 6974 80000
rect 9678 79200 9734 80000
rect 12438 79200 12494 80000
rect 15198 79200 15254 80000
rect 17958 79200 18014 80000
rect 20718 79200 20774 80000
rect 23478 79200 23534 80000
rect 26238 79200 26294 80000
rect 28998 79200 29054 80000
rect 31758 79200 31814 80000
rect 34518 79200 34574 80000
rect 37278 79200 37334 80000
rect 40038 79200 40094 80000
rect 42798 79200 42854 80000
rect 45558 79200 45614 80000
rect 48318 79200 48374 80000
rect 51078 79200 51134 80000
rect 53838 79200 53894 80000
rect 56598 79200 56654 80000
rect 59358 79200 59414 80000
rect 62118 79200 62174 80000
rect 64878 79200 64934 80000
rect 67638 79200 67694 80000
rect 70398 79200 70454 80000
rect 73158 79200 73214 80000
rect 75918 79200 75974 80000
rect 78678 79200 78734 80000
rect 1582 0 1638 800
rect 4710 0 4766 800
rect 7930 0 7986 800
rect 11150 0 11206 800
rect 14370 0 14426 800
rect 17590 0 17646 800
rect 20718 0 20774 800
rect 23938 0 23994 800
rect 27158 0 27214 800
rect 30378 0 30434 800
rect 33598 0 33654 800
rect 36726 0 36782 800
rect 39946 0 40002 800
rect 43166 0 43222 800
rect 46386 0 46442 800
rect 49606 0 49662 800
rect 52734 0 52790 800
rect 55954 0 56010 800
rect 59174 0 59230 800
rect 62394 0 62450 800
rect 65614 0 65670 800
rect 68742 0 68798 800
rect 71962 0 72018 800
rect 75182 0 75238 800
rect 78402 0 78458 800
<< obsm2 >>
rect 1510 79144 4102 79200
rect 4270 79144 6862 79200
rect 7030 79144 9622 79200
rect 9790 79144 12382 79200
rect 12550 79144 15142 79200
rect 15310 79144 17902 79200
rect 18070 79144 20662 79200
rect 20830 79144 23422 79200
rect 23590 79144 26182 79200
rect 26350 79144 28942 79200
rect 29110 79144 31702 79200
rect 31870 79144 34462 79200
rect 34630 79144 37222 79200
rect 37390 79144 39982 79200
rect 40150 79144 42742 79200
rect 42910 79144 45502 79200
rect 45670 79144 48262 79200
rect 48430 79144 51022 79200
rect 51190 79144 53782 79200
rect 53950 79144 56542 79200
rect 56710 79144 59302 79200
rect 59470 79144 62062 79200
rect 62230 79144 64822 79200
rect 64990 79144 67582 79200
rect 67750 79144 70342 79200
rect 70510 79144 73102 79200
rect 73270 79144 75862 79200
rect 76030 79144 78622 79200
rect 1398 856 78732 79144
rect 1398 800 1526 856
rect 1694 800 4654 856
rect 4822 800 7874 856
rect 8042 800 11094 856
rect 11262 800 14314 856
rect 14482 800 17534 856
rect 17702 800 20662 856
rect 20830 800 23882 856
rect 24050 800 27102 856
rect 27270 800 30322 856
rect 30490 800 33542 856
rect 33710 800 36670 856
rect 36838 800 39890 856
rect 40058 800 43110 856
rect 43278 800 46330 856
rect 46498 800 49550 856
rect 49718 800 52678 856
rect 52846 800 55898 856
rect 56066 800 59118 856
rect 59286 800 62338 856
rect 62506 800 65558 856
rect 65726 800 68686 856
rect 68854 800 71906 856
rect 72074 800 75126 856
rect 75294 800 78346 856
rect 78514 800 78732 856
<< metal3 >>
rect 0 78072 800 78192
rect 79200 77800 80000 77920
rect 0 74400 800 74520
rect 79200 73584 80000 73704
rect 0 70728 800 70848
rect 79200 69368 80000 69488
rect 0 67192 800 67312
rect 79200 65152 80000 65272
rect 0 63520 800 63640
rect 79200 60936 80000 61056
rect 0 59848 800 59968
rect 79200 56720 80000 56840
rect 0 56176 800 56296
rect 0 52640 800 52760
rect 79200 52504 80000 52624
rect 0 48968 800 49088
rect 79200 48288 80000 48408
rect 0 45296 800 45416
rect 79200 44072 80000 44192
rect 0 41760 800 41880
rect 79200 39856 80000 39976
rect 0 38088 800 38208
rect 79200 35640 80000 35760
rect 0 34416 800 34536
rect 79200 31424 80000 31544
rect 0 30744 800 30864
rect 0 27208 800 27328
rect 79200 27208 80000 27328
rect 0 23536 800 23656
rect 79200 22992 80000 23112
rect 0 19864 800 19984
rect 79200 18776 80000 18896
rect 0 16192 800 16312
rect 79200 14560 80000 14680
rect 0 12656 800 12776
rect 79200 10344 80000 10464
rect 0 8984 800 9104
rect 79200 6128 80000 6248
rect 0 5312 800 5432
rect 79200 2048 80000 2168
rect 0 1776 800 1896
<< obsm3 >>
rect 880 78000 79200 78165
rect 880 77992 79120 78000
rect 800 77720 79120 77992
rect 800 74600 79200 77720
rect 880 74320 79200 74600
rect 800 73784 79200 74320
rect 800 73504 79120 73784
rect 800 70928 79200 73504
rect 880 70648 79200 70928
rect 800 69568 79200 70648
rect 800 69288 79120 69568
rect 800 67392 79200 69288
rect 880 67112 79200 67392
rect 800 65352 79200 67112
rect 800 65072 79120 65352
rect 800 63720 79200 65072
rect 880 63440 79200 63720
rect 800 61136 79200 63440
rect 800 60856 79120 61136
rect 800 60048 79200 60856
rect 880 59768 79200 60048
rect 800 56920 79200 59768
rect 800 56640 79120 56920
rect 800 56376 79200 56640
rect 880 56096 79200 56376
rect 800 52840 79200 56096
rect 880 52704 79200 52840
rect 880 52560 79120 52704
rect 800 52424 79120 52560
rect 800 49168 79200 52424
rect 880 48888 79200 49168
rect 800 48488 79200 48888
rect 800 48208 79120 48488
rect 800 45496 79200 48208
rect 880 45216 79200 45496
rect 800 44272 79200 45216
rect 800 43992 79120 44272
rect 800 41960 79200 43992
rect 880 41680 79200 41960
rect 800 40056 79200 41680
rect 800 39776 79120 40056
rect 800 38288 79200 39776
rect 880 38008 79200 38288
rect 800 35840 79200 38008
rect 800 35560 79120 35840
rect 800 34616 79200 35560
rect 880 34336 79200 34616
rect 800 31624 79200 34336
rect 800 31344 79120 31624
rect 800 30944 79200 31344
rect 880 30664 79200 30944
rect 800 27408 79200 30664
rect 880 27128 79120 27408
rect 800 23736 79200 27128
rect 880 23456 79200 23736
rect 800 23192 79200 23456
rect 800 22912 79120 23192
rect 800 20064 79200 22912
rect 880 19784 79200 20064
rect 800 18976 79200 19784
rect 800 18696 79120 18976
rect 800 16392 79200 18696
rect 880 16112 79200 16392
rect 800 14760 79200 16112
rect 800 14480 79120 14760
rect 800 12856 79200 14480
rect 880 12576 79200 12856
rect 800 10544 79200 12576
rect 800 10264 79120 10544
rect 800 9184 79200 10264
rect 880 8904 79200 9184
rect 800 6328 79200 8904
rect 800 6048 79120 6328
rect 800 5512 79200 6048
rect 880 5232 79200 5512
rect 800 2248 79200 5232
rect 800 1976 79120 2248
rect 880 1968 79120 1976
rect 880 1803 79200 1968
<< metal4 >>
rect 4208 2128 4528 77840
rect 19568 2128 19888 77840
rect 34928 2128 35248 77840
rect 50288 2128 50608 77840
rect 65648 2128 65968 77840
<< obsm4 >>
rect 15515 2347 19488 77349
rect 19968 2347 34848 77349
rect 35328 2347 50208 77349
rect 50688 2347 65568 77349
rect 66048 2347 67837 77349
<< labels >>
rlabel metal2 s 1582 0 1638 800 6 clock
port 1 nsew signal input
rlabel metal2 s 7930 0 7986 800 6 io_ba_match
port 2 nsew signal input
rlabel metal3 s 0 1776 800 1896 6 io_motor_irq
port 3 nsew signal output
rlabel metal2 s 1398 79200 1454 80000 6 io_pwm_high
port 4 nsew signal output
rlabel metal2 s 4158 79200 4214 80000 6 io_pwm_low
port 5 nsew signal output
rlabel metal2 s 6918 79200 6974 80000 6 io_qei_ch_a
port 6 nsew signal input
rlabel metal3 s 79200 2048 80000 2168 6 io_qei_ch_b
port 7 nsew signal input
rlabel metal2 s 9678 79200 9734 80000 6 io_wbs_ack_o
port 8 nsew signal output
rlabel metal2 s 15198 79200 15254 80000 6 io_wbs_data_o[0]
port 9 nsew signal output
rlabel metal2 s 39946 0 40002 800 6 io_wbs_data_o[10]
port 10 nsew signal output
rlabel metal2 s 48318 79200 48374 80000 6 io_wbs_data_o[11]
port 11 nsew signal output
rlabel metal2 s 43166 0 43222 800 6 io_wbs_data_o[12]
port 12 nsew signal output
rlabel metal3 s 79200 39856 80000 39976 6 io_wbs_data_o[13]
port 13 nsew signal output
rlabel metal2 s 49606 0 49662 800 6 io_wbs_data_o[14]
port 14 nsew signal output
rlabel metal2 s 55954 0 56010 800 6 io_wbs_data_o[15]
port 15 nsew signal output
rlabel metal3 s 79200 52504 80000 52624 6 io_wbs_data_o[16]
port 16 nsew signal output
rlabel metal3 s 79200 56720 80000 56840 6 io_wbs_data_o[17]
port 17 nsew signal output
rlabel metal2 s 62394 0 62450 800 6 io_wbs_data_o[18]
port 18 nsew signal output
rlabel metal3 s 0 56176 800 56296 6 io_wbs_data_o[19]
port 19 nsew signal output
rlabel metal2 s 20718 79200 20774 80000 6 io_wbs_data_o[1]
port 20 nsew signal output
rlabel metal2 s 56598 79200 56654 80000 6 io_wbs_data_o[20]
port 21 nsew signal output
rlabel metal3 s 0 63520 800 63640 6 io_wbs_data_o[21]
port 22 nsew signal output
rlabel metal2 s 65614 0 65670 800 6 io_wbs_data_o[22]
port 23 nsew signal output
rlabel metal3 s 0 67192 800 67312 6 io_wbs_data_o[23]
port 24 nsew signal output
rlabel metal2 s 68742 0 68798 800 6 io_wbs_data_o[24]
port 25 nsew signal output
rlabel metal2 s 71962 0 72018 800 6 io_wbs_data_o[25]
port 26 nsew signal output
rlabel metal2 s 70398 79200 70454 80000 6 io_wbs_data_o[26]
port 27 nsew signal output
rlabel metal2 s 73158 79200 73214 80000 6 io_wbs_data_o[27]
port 28 nsew signal output
rlabel metal2 s 75182 0 75238 800 6 io_wbs_data_o[28]
port 29 nsew signal output
rlabel metal2 s 75918 79200 75974 80000 6 io_wbs_data_o[29]
port 30 nsew signal output
rlabel metal3 s 0 8984 800 9104 6 io_wbs_data_o[2]
port 31 nsew signal output
rlabel metal2 s 78678 79200 78734 80000 6 io_wbs_data_o[30]
port 32 nsew signal output
rlabel metal3 s 79200 77800 80000 77920 6 io_wbs_data_o[31]
port 33 nsew signal output
rlabel metal2 s 23478 79200 23534 80000 6 io_wbs_data_o[3]
port 34 nsew signal output
rlabel metal2 s 23938 0 23994 800 6 io_wbs_data_o[4]
port 35 nsew signal output
rlabel metal2 s 31758 79200 31814 80000 6 io_wbs_data_o[5]
port 36 nsew signal output
rlabel metal3 s 79200 18776 80000 18896 6 io_wbs_data_o[6]
port 37 nsew signal output
rlabel metal2 s 37278 79200 37334 80000 6 io_wbs_data_o[7]
port 38 nsew signal output
rlabel metal2 s 30378 0 30434 800 6 io_wbs_data_o[8]
port 39 nsew signal output
rlabel metal2 s 36726 0 36782 800 6 io_wbs_data_o[9]
port 40 nsew signal output
rlabel metal2 s 14370 0 14426 800 6 io_wbs_m2s_addr[0]
port 41 nsew signal input
rlabel metal3 s 79200 27208 80000 27328 6 io_wbs_m2s_addr[10]
port 42 nsew signal input
rlabel metal3 s 79200 31424 80000 31544 6 io_wbs_m2s_addr[11]
port 43 nsew signal input
rlabel metal2 s 46386 0 46442 800 6 io_wbs_m2s_addr[12]
port 44 nsew signal input
rlabel metal3 s 79200 44072 80000 44192 6 io_wbs_m2s_addr[13]
port 45 nsew signal input
rlabel metal3 s 0 45296 800 45416 6 io_wbs_m2s_addr[14]
port 46 nsew signal input
rlabel metal3 s 79200 48288 80000 48408 6 io_wbs_m2s_addr[15]
port 47 nsew signal input
rlabel metal3 s 0 5312 800 5432 6 io_wbs_m2s_addr[1]
port 48 nsew signal input
rlabel metal3 s 0 12656 800 12776 6 io_wbs_m2s_addr[2]
port 49 nsew signal input
rlabel metal2 s 26238 79200 26294 80000 6 io_wbs_m2s_addr[3]
port 50 nsew signal input
rlabel metal3 s 79200 14560 80000 14680 6 io_wbs_m2s_addr[4]
port 51 nsew signal input
rlabel metal2 s 34518 79200 34574 80000 6 io_wbs_m2s_addr[5]
port 52 nsew signal input
rlabel metal3 s 0 27208 800 27328 6 io_wbs_m2s_addr[6]
port 53 nsew signal input
rlabel metal3 s 0 34416 800 34536 6 io_wbs_m2s_addr[7]
port 54 nsew signal input
rlabel metal2 s 33598 0 33654 800 6 io_wbs_m2s_addr[8]
port 55 nsew signal input
rlabel metal3 s 79200 22992 80000 23112 6 io_wbs_m2s_addr[9]
port 56 nsew signal input
rlabel metal2 s 17590 0 17646 800 6 io_wbs_m2s_data[0]
port 57 nsew signal input
rlabel metal2 s 45558 79200 45614 80000 6 io_wbs_m2s_data[10]
port 58 nsew signal input
rlabel metal3 s 79200 35640 80000 35760 6 io_wbs_m2s_data[11]
port 59 nsew signal input
rlabel metal2 s 51078 79200 51134 80000 6 io_wbs_m2s_data[12]
port 60 nsew signal input
rlabel metal3 s 0 41760 800 41880 6 io_wbs_m2s_data[13]
port 61 nsew signal input
rlabel metal2 s 52734 0 52790 800 6 io_wbs_m2s_data[14]
port 62 nsew signal input
rlabel metal2 s 59174 0 59230 800 6 io_wbs_m2s_data[15]
port 63 nsew signal input
rlabel metal3 s 0 48968 800 49088 6 io_wbs_m2s_data[16]
port 64 nsew signal input
rlabel metal2 s 53838 79200 53894 80000 6 io_wbs_m2s_data[17]
port 65 nsew signal input
rlabel metal3 s 0 52640 800 52760 6 io_wbs_m2s_data[18]
port 66 nsew signal input
rlabel metal3 s 0 59848 800 59968 6 io_wbs_m2s_data[19]
port 67 nsew signal input
rlabel metal3 s 79200 6128 80000 6248 6 io_wbs_m2s_data[1]
port 68 nsew signal input
rlabel metal3 s 79200 60936 80000 61056 6 io_wbs_m2s_data[20]
port 69 nsew signal input
rlabel metal2 s 59358 79200 59414 80000 6 io_wbs_m2s_data[21]
port 70 nsew signal input
rlabel metal2 s 62118 79200 62174 80000 6 io_wbs_m2s_data[22]
port 71 nsew signal input
rlabel metal3 s 79200 65152 80000 65272 6 io_wbs_m2s_data[23]
port 72 nsew signal input
rlabel metal2 s 64878 79200 64934 80000 6 io_wbs_m2s_data[24]
port 73 nsew signal input
rlabel metal2 s 67638 79200 67694 80000 6 io_wbs_m2s_data[25]
port 74 nsew signal input
rlabel metal3 s 79200 69368 80000 69488 6 io_wbs_m2s_data[26]
port 75 nsew signal input
rlabel metal3 s 0 70728 800 70848 6 io_wbs_m2s_data[27]
port 76 nsew signal input
rlabel metal2 s 78402 0 78458 800 6 io_wbs_m2s_data[28]
port 77 nsew signal input
rlabel metal3 s 0 74400 800 74520 6 io_wbs_m2s_data[29]
port 78 nsew signal input
rlabel metal3 s 0 16192 800 16312 6 io_wbs_m2s_data[2]
port 79 nsew signal input
rlabel metal3 s 79200 73584 80000 73704 6 io_wbs_m2s_data[30]
port 80 nsew signal input
rlabel metal3 s 0 78072 800 78192 6 io_wbs_m2s_data[31]
port 81 nsew signal input
rlabel metal2 s 28998 79200 29054 80000 6 io_wbs_m2s_data[3]
port 82 nsew signal input
rlabel metal3 s 0 23536 800 23656 6 io_wbs_m2s_data[4]
port 83 nsew signal input
rlabel metal2 s 27158 0 27214 800 6 io_wbs_m2s_data[5]
port 84 nsew signal input
rlabel metal3 s 0 30744 800 30864 6 io_wbs_m2s_data[6]
port 85 nsew signal input
rlabel metal2 s 40038 79200 40094 80000 6 io_wbs_m2s_data[7]
port 86 nsew signal input
rlabel metal2 s 42798 79200 42854 80000 6 io_wbs_m2s_data[8]
port 87 nsew signal input
rlabel metal3 s 0 38088 800 38208 6 io_wbs_m2s_data[9]
port 88 nsew signal input
rlabel metal2 s 17958 79200 18014 80000 6 io_wbs_m2s_sel[0]
port 89 nsew signal input
rlabel metal3 s 79200 10344 80000 10464 6 io_wbs_m2s_sel[1]
port 90 nsew signal input
rlabel metal3 s 0 19864 800 19984 6 io_wbs_m2s_sel[2]
port 91 nsew signal input
rlabel metal2 s 20718 0 20774 800 6 io_wbs_m2s_sel[3]
port 92 nsew signal input
rlabel metal2 s 11150 0 11206 800 6 io_wbs_m2s_stb
port 93 nsew signal input
rlabel metal2 s 12438 79200 12494 80000 6 io_wbs_m2s_we
port 94 nsew signal input
rlabel metal2 s 4710 0 4766 800 6 reset
port 95 nsew signal input
rlabel metal4 s 4208 2128 4528 77840 6 vccd1
port 96 nsew power input
rlabel metal4 s 34928 2128 35248 77840 6 vccd1
port 96 nsew power input
rlabel metal4 s 65648 2128 65968 77840 6 vccd1
port 96 nsew power input
rlabel metal4 s 19568 2128 19888 77840 6 vssd1
port 97 nsew ground input
rlabel metal4 s 50288 2128 50608 77840 6 vssd1
port 97 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 80000 80000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 16647140
string GDS_FILE /home/em/mpw/UETRV-ECORE/openlane/Motor_Top/runs/Motor_Top/results/finishing/Motor_Top.magic.gds
string GDS_START 1021908
<< end >>

