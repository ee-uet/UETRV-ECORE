magic
tech sky130A
magscale 1 2
timestamp 1647682248
<< viali >>
rect 4169 33609 4203 33643
rect 6745 33609 6779 33643
rect 9873 33609 9907 33643
rect 16957 33609 16991 33643
rect 18245 33609 18279 33643
rect 23029 33609 23063 33643
rect 23949 33609 23983 33643
rect 26065 33609 26099 33643
rect 26525 33609 26559 33643
rect 28181 33609 28215 33643
rect 29101 33609 29135 33643
rect 29929 33609 29963 33643
rect 31769 33609 31803 33643
rect 2789 33541 2823 33575
rect 3249 33541 3283 33575
rect 17417 33541 17451 33575
rect 32505 33541 32539 33575
rect 2237 33473 2271 33507
rect 2973 33473 3007 33507
rect 3985 33473 4019 33507
rect 4629 33473 4663 33507
rect 5733 33473 5767 33507
rect 6561 33473 6595 33507
rect 7941 33473 7975 33507
rect 8401 33473 8435 33507
rect 9229 33473 9263 33507
rect 10057 33473 10091 33507
rect 10885 33473 10919 33507
rect 11713 33473 11747 33507
rect 12173 33473 12207 33507
rect 13737 33473 13771 33507
rect 14381 33473 14415 33507
rect 14657 33473 14691 33507
rect 15117 33473 15151 33507
rect 16037 33473 16071 33507
rect 17141 33473 17175 33507
rect 18429 33473 18463 33507
rect 18889 33473 18923 33507
rect 19441 33473 19475 33507
rect 20637 33473 20671 33507
rect 20913 33473 20947 33507
rect 21833 33473 21867 33507
rect 22293 33473 22327 33507
rect 23489 33473 23523 33507
rect 24409 33473 24443 33507
rect 25605 33473 25639 33507
rect 25881 33473 25915 33507
rect 26985 33473 27019 33507
rect 28457 33473 28491 33507
rect 28917 33473 28951 33507
rect 29745 33473 29779 33507
rect 30389 33473 30423 33507
rect 33149 33473 33183 33507
rect 1961 33405 1995 33439
rect 4905 33405 4939 33439
rect 11161 33405 11195 33439
rect 16313 33405 16347 33439
rect 19717 33405 19751 33439
rect 24685 33405 24719 33439
rect 27261 33405 27295 33439
rect 30665 33405 30699 33439
rect 33517 33405 33551 33439
rect 33793 33405 33827 33439
rect 5917 33337 5951 33371
rect 14197 33337 14231 33371
rect 14841 33337 14875 33371
rect 23305 33337 23339 33371
rect 32321 33337 32355 33371
rect 32965 33337 32999 33371
rect 8033 33269 8067 33303
rect 9321 33269 9355 33303
rect 11897 33269 11931 33303
rect 22017 33269 22051 33303
rect 28641 33269 28675 33303
rect 2789 33065 2823 33099
rect 4537 33065 4571 33099
rect 5549 33065 5583 33099
rect 6009 33065 6043 33099
rect 8493 33065 8527 33099
rect 10793 33065 10827 33099
rect 11529 33065 11563 33099
rect 14657 33065 14691 33099
rect 16405 33065 16439 33099
rect 16957 33065 16991 33099
rect 19441 33065 19475 33099
rect 21557 33065 21591 33099
rect 24685 33065 24719 33099
rect 25421 33065 25455 33099
rect 27261 33065 27295 33099
rect 30297 33065 30331 33099
rect 30757 33065 30791 33099
rect 32505 33065 32539 33099
rect 33149 33065 33183 33099
rect 33701 33065 33735 33099
rect 3157 32997 3191 33031
rect 17417 32997 17451 33031
rect 22109 32997 22143 33031
rect 27721 32997 27755 33031
rect 14933 32929 14967 32963
rect 31033 32929 31067 32963
rect 1685 32861 1719 32895
rect 2237 32861 2271 32895
rect 3341 32861 3375 32895
rect 6193 32861 6227 32895
rect 9321 32861 9355 32895
rect 9597 32861 9631 32895
rect 11069 32861 11103 32895
rect 15209 32861 15243 32895
rect 16221 32861 16255 32895
rect 16773 32861 16807 32895
rect 17601 32861 17635 32895
rect 18061 32861 18095 32895
rect 19257 32861 19291 32895
rect 21925 32861 21959 32895
rect 24869 32861 24903 32895
rect 25237 32861 25271 32895
rect 27445 32861 27479 32895
rect 27905 32861 27939 32895
rect 31309 32861 31343 32895
rect 32321 32861 32355 32895
rect 32965 32861 32999 32895
rect 33517 32861 33551 32895
rect 34253 32861 34287 32895
rect 1869 32793 1903 32827
rect 17877 32793 17911 32827
rect 18521 32793 18555 32827
rect 2329 32725 2363 32759
rect 6469 32725 6503 32759
rect 9137 32725 9171 32759
rect 11253 32725 11287 32759
rect 18613 32725 18647 32759
rect 28733 32725 28767 32759
rect 34161 32725 34195 32759
rect 2605 32521 2639 32555
rect 15577 32521 15611 32555
rect 32781 32521 32815 32555
rect 33057 32521 33091 32555
rect 33701 32521 33735 32555
rect 3065 32453 3099 32487
rect 17877 32453 17911 32487
rect 18061 32453 18095 32487
rect 2789 32385 2823 32419
rect 15393 32385 15427 32419
rect 18521 32385 18555 32419
rect 18981 32385 19015 32419
rect 33241 32385 33275 32419
rect 33517 32385 33551 32419
rect 34069 32385 34103 32419
rect 1409 32317 1443 32351
rect 1685 32317 1719 32351
rect 32413 32317 32447 32351
rect 18705 32249 18739 32283
rect 31769 32181 31803 32215
rect 34253 32181 34287 32215
rect 2053 31977 2087 32011
rect 32965 31977 32999 32011
rect 33333 31977 33367 32011
rect 34253 31977 34287 32011
rect 2605 31909 2639 31943
rect 33793 31909 33827 31943
rect 1685 31773 1719 31807
rect 2237 31773 2271 31807
rect 2973 31773 3007 31807
rect 32597 31773 32631 31807
rect 33609 31773 33643 31807
rect 34069 31773 34103 31807
rect 1501 31637 1535 31671
rect 1409 31433 1443 31467
rect 17877 31365 17911 31399
rect 33885 31297 33919 31331
rect 34345 31297 34379 31331
rect 17969 31093 18003 31127
rect 33425 31093 33459 31127
rect 34161 31093 34195 31127
rect 34069 30753 34103 30787
rect 1685 30685 1719 30719
rect 34345 30685 34379 30719
rect 1501 30549 1535 30583
rect 2053 30549 2087 30583
rect 33885 30345 33919 30379
rect 1961 30209 1995 30243
rect 33517 30209 33551 30243
rect 34345 30209 34379 30243
rect 2237 30141 2271 30175
rect 34161 30005 34195 30039
rect 1961 29801 1995 29835
rect 34161 29801 34195 29835
rect 1685 29597 1719 29631
rect 33885 29597 33919 29631
rect 34345 29597 34379 29631
rect 1501 29461 1535 29495
rect 2421 29461 2455 29495
rect 1685 29121 1719 29155
rect 2145 29121 2179 29155
rect 33609 29121 33643 29155
rect 34069 29121 34103 29155
rect 1869 28985 1903 29019
rect 34253 28985 34287 29019
rect 33793 28917 33827 28951
rect 33977 28713 34011 28747
rect 20269 28169 20303 28203
rect 1685 28033 1719 28067
rect 30941 28033 30975 28067
rect 34069 28033 34103 28067
rect 1501 27897 1535 27931
rect 34253 27897 34287 27931
rect 2053 27829 2087 27863
rect 31125 27829 31159 27863
rect 19901 27557 19935 27591
rect 20913 27489 20947 27523
rect 19625 27421 19659 27455
rect 19809 27421 19843 27455
rect 19993 27421 20027 27455
rect 20085 27421 20119 27455
rect 20453 27421 20487 27455
rect 20637 27421 20671 27455
rect 21281 27421 21315 27455
rect 19257 27285 19291 27319
rect 20545 27285 20579 27319
rect 21649 27285 21683 27319
rect 18613 27081 18647 27115
rect 19625 27081 19659 27115
rect 21189 27081 21223 27115
rect 17969 26945 18003 26979
rect 19533 26945 19567 26979
rect 19901 26945 19935 26979
rect 20085 26945 20119 26979
rect 20729 26945 20763 26979
rect 21189 26945 21223 26979
rect 21373 26945 21407 26979
rect 33793 26945 33827 26979
rect 34253 26945 34287 26979
rect 20637 26877 20671 26911
rect 21833 26877 21867 26911
rect 17785 26809 17819 26843
rect 18981 26741 19015 26775
rect 20361 26741 20395 26775
rect 22293 26741 22327 26775
rect 34161 26741 34195 26775
rect 18245 26537 18279 26571
rect 21281 26537 21315 26571
rect 21465 26537 21499 26571
rect 1593 26469 1627 26503
rect 18797 26469 18831 26503
rect 34161 26469 34195 26503
rect 19625 26401 19659 26435
rect 20545 26401 20579 26435
rect 21925 26401 21959 26435
rect 1409 26333 1443 26367
rect 1869 26333 1903 26367
rect 18705 26333 18739 26367
rect 19809 26333 19843 26367
rect 19993 26333 20027 26367
rect 20085 26333 20119 26367
rect 20269 26333 20303 26367
rect 20729 26333 20763 26367
rect 21005 26333 21039 26367
rect 33885 26333 33919 26367
rect 34345 26333 34379 26367
rect 19901 26265 19935 26299
rect 21649 26265 21683 26299
rect 20913 26197 20947 26231
rect 21449 26197 21483 26231
rect 18981 25993 19015 26027
rect 19625 25993 19659 26027
rect 20361 25993 20395 26027
rect 17877 25925 17911 25959
rect 19257 25925 19291 25959
rect 19473 25925 19507 25959
rect 18613 25857 18647 25891
rect 20085 25857 20119 25891
rect 20453 25857 20487 25891
rect 21281 25857 21315 25891
rect 19901 25789 19935 25823
rect 20821 25789 20855 25823
rect 17969 25653 18003 25687
rect 19441 25653 19475 25687
rect 21005 25653 21039 25687
rect 21833 25653 21867 25687
rect 19257 25449 19291 25483
rect 19901 25449 19935 25483
rect 20085 25449 20119 25483
rect 6285 25245 6319 25279
rect 19441 25245 19475 25279
rect 20545 25245 20579 25279
rect 20729 25245 20763 25279
rect 34069 25245 34103 25279
rect 20053 25177 20087 25211
rect 20269 25177 20303 25211
rect 6101 25109 6135 25143
rect 20637 25109 20671 25143
rect 21005 25109 21039 25143
rect 34253 25109 34287 25143
rect 19809 24905 19843 24939
rect 1685 24769 1719 24803
rect 34069 24769 34103 24803
rect 1501 24565 1535 24599
rect 2053 24565 2087 24599
rect 20453 24565 20487 24599
rect 34253 24565 34287 24599
rect 1685 24157 1719 24191
rect 2053 24089 2087 24123
rect 33977 24089 34011 24123
rect 34161 24089 34195 24123
rect 1501 24021 1535 24055
rect 33609 24021 33643 24055
rect 33793 23749 33827 23783
rect 34253 23749 34287 23783
rect 1685 23681 1719 23715
rect 34069 23545 34103 23579
rect 1501 23477 1535 23511
rect 33701 23273 33735 23307
rect 34253 23205 34287 23239
rect 34069 23069 34103 23103
rect 1685 22593 1719 22627
rect 18061 22593 18095 22627
rect 34069 22593 34103 22627
rect 34345 22525 34379 22559
rect 1501 22457 1535 22491
rect 17877 22457 17911 22491
rect 33977 22185 34011 22219
rect 34345 21845 34379 21879
rect 1685 21505 1719 21539
rect 34069 21505 34103 21539
rect 34345 21437 34379 21471
rect 1501 21301 1535 21335
rect 33241 20893 33275 20927
rect 33517 20893 33551 20927
rect 33793 20893 33827 20927
rect 17969 20825 18003 20859
rect 17877 20757 17911 20791
rect 33977 20553 34011 20587
rect 34161 20417 34195 20451
rect 1409 20213 1443 20247
rect 34161 20009 34195 20043
rect 1409 19805 1443 19839
rect 1685 19805 1719 19839
rect 33885 19805 33919 19839
rect 34345 19805 34379 19839
rect 1593 19465 1627 19499
rect 34161 19465 34195 19499
rect 17969 19397 18003 19431
rect 1409 19329 1443 19363
rect 1961 19329 1995 19363
rect 18521 19329 18555 19363
rect 18981 19329 19015 19363
rect 33885 19329 33919 19363
rect 34345 19329 34379 19363
rect 18705 19193 18739 19227
rect 17233 19125 17267 19159
rect 18061 19125 18095 19159
rect 29745 18853 29779 18887
rect 17049 18785 17083 18819
rect 1685 18717 1719 18751
rect 2145 18717 2179 18751
rect 2421 18717 2455 18751
rect 17417 18717 17451 18751
rect 17969 18717 18003 18751
rect 18613 18717 18647 18751
rect 20729 18717 20763 18751
rect 21189 18717 21223 18751
rect 29561 18717 29595 18751
rect 33885 18717 33919 18751
rect 34345 18717 34379 18751
rect 18153 18649 18187 18683
rect 23213 18649 23247 18683
rect 23397 18649 23431 18683
rect 1501 18581 1535 18615
rect 1961 18581 1995 18615
rect 17509 18581 17543 18615
rect 18521 18581 18555 18615
rect 19349 18581 19383 18615
rect 20821 18581 20855 18615
rect 34161 18581 34195 18615
rect 2237 18377 2271 18411
rect 3525 18377 3559 18411
rect 7113 18377 7147 18411
rect 12909 18377 12943 18411
rect 16221 18377 16255 18411
rect 17969 18377 18003 18411
rect 29193 18377 29227 18411
rect 29929 18377 29963 18411
rect 1777 18309 1811 18343
rect 3065 18309 3099 18343
rect 5549 18309 5583 18343
rect 6561 18309 6595 18343
rect 17325 18309 17359 18343
rect 18521 18309 18555 18343
rect 24501 18309 24535 18343
rect 27629 18309 27663 18343
rect 29561 18309 29595 18343
rect 31217 18309 31251 18343
rect 32505 18309 32539 18343
rect 2421 18241 2455 18275
rect 3617 18241 3651 18275
rect 6745 18241 6779 18275
rect 7297 18241 7331 18275
rect 13093 18241 13127 18275
rect 15853 18241 15887 18275
rect 16773 18241 16807 18275
rect 17877 18241 17911 18275
rect 18981 18241 19015 18275
rect 19533 18241 19567 18275
rect 27445 18241 27479 18275
rect 29377 18241 29411 18275
rect 30021 18241 30055 18275
rect 33609 18241 33643 18275
rect 34069 18241 34103 18275
rect 19993 18173 20027 18207
rect 5733 18105 5767 18139
rect 15669 18105 15703 18139
rect 16957 18105 16991 18139
rect 17509 18105 17543 18139
rect 19717 18105 19751 18139
rect 24685 18105 24719 18139
rect 32321 18105 32355 18139
rect 1869 18037 1903 18071
rect 2973 18037 3007 18071
rect 18429 18037 18463 18071
rect 19073 18037 19107 18071
rect 30389 18037 30423 18071
rect 31309 18037 31343 18071
rect 33793 18037 33827 18071
rect 34253 18037 34287 18071
rect 2605 17833 2639 17867
rect 16037 17833 16071 17867
rect 16681 17833 16715 17867
rect 17049 17833 17083 17867
rect 18521 17833 18555 17867
rect 1777 17629 1811 17663
rect 17417 17629 17451 17663
rect 17969 17629 18003 17663
rect 19717 17629 19751 17663
rect 29837 17629 29871 17663
rect 30297 17629 30331 17663
rect 2513 17561 2547 17595
rect 17601 17561 17635 17595
rect 18613 17561 18647 17595
rect 19533 17561 19567 17595
rect 30021 17561 30055 17595
rect 1869 17493 1903 17527
rect 18061 17493 18095 17527
rect 17417 17289 17451 17323
rect 17969 17289 18003 17323
rect 30021 17289 30055 17323
rect 33793 17289 33827 17323
rect 18337 17221 18371 17255
rect 18521 17221 18555 17255
rect 1685 17153 1719 17187
rect 17877 17153 17911 17187
rect 29837 17153 29871 17187
rect 33609 17153 33643 17187
rect 34069 17153 34103 17187
rect 18981 17085 19015 17119
rect 1501 17017 1535 17051
rect 34253 17017 34287 17051
rect 17693 16745 17727 16779
rect 34345 16405 34379 16439
rect 1685 16065 1719 16099
rect 34069 15997 34103 16031
rect 34345 15997 34379 16031
rect 1501 15861 1535 15895
rect 1593 15657 1627 15691
rect 1409 15453 1443 15487
rect 1869 15453 1903 15487
rect 34069 15453 34103 15487
rect 34253 15317 34287 15351
rect 18521 15113 18555 15147
rect 33977 15113 34011 15147
rect 18061 15045 18095 15079
rect 18613 14977 18647 15011
rect 34161 14977 34195 15011
rect 17877 14841 17911 14875
rect 18981 14773 19015 14807
rect 34161 14569 34195 14603
rect 1685 14365 1719 14399
rect 33517 14365 33551 14399
rect 34345 14365 34379 14399
rect 1501 14229 1535 14263
rect 33885 14229 33919 14263
rect 34069 13889 34103 13923
rect 34345 13821 34379 13855
rect 34069 13277 34103 13311
rect 1685 13209 1719 13243
rect 1869 13209 1903 13243
rect 2145 13141 2179 13175
rect 33701 13141 33735 13175
rect 34253 13141 34287 13175
rect 1685 12801 1719 12835
rect 33701 12801 33735 12835
rect 34069 12801 34103 12835
rect 1501 12597 1535 12631
rect 2053 12597 2087 12631
rect 34253 12597 34287 12631
rect 17969 11713 18003 11747
rect 34069 11713 34103 11747
rect 1409 11645 1443 11679
rect 1685 11645 1719 11679
rect 18153 11645 18187 11679
rect 34253 11577 34287 11611
rect 1409 11305 1443 11339
rect 1593 10761 1627 10795
rect 1409 10625 1443 10659
rect 1869 10625 1903 10659
rect 34161 10217 34195 10251
rect 33885 10013 33919 10047
rect 34345 10013 34379 10047
rect 17417 9945 17451 9979
rect 17509 9877 17543 9911
rect 18061 9537 18095 9571
rect 17877 9401 17911 9435
rect 18521 9333 18555 9367
rect 1685 8925 1719 8959
rect 33701 8925 33735 8959
rect 34069 8925 34103 8959
rect 2053 8857 2087 8891
rect 1501 8789 1535 8823
rect 34253 8789 34287 8823
rect 33793 8449 33827 8483
rect 34253 8449 34287 8483
rect 34069 8313 34103 8347
rect 1685 7837 1719 7871
rect 34069 7837 34103 7871
rect 1501 7701 1535 7735
rect 34253 7701 34287 7735
rect 1685 7361 1719 7395
rect 34069 7361 34103 7395
rect 1501 7157 1535 7191
rect 2053 7157 2087 7191
rect 34253 7157 34287 7191
rect 1685 6273 1719 6307
rect 33793 6273 33827 6307
rect 34253 6273 34287 6307
rect 1501 6137 1535 6171
rect 34069 6137 34103 6171
rect 34345 5525 34379 5559
rect 10977 5321 11011 5355
rect 1685 5185 1719 5219
rect 11161 5185 11195 5219
rect 34069 5117 34103 5151
rect 34345 5117 34379 5151
rect 1501 4981 1535 5015
rect 17877 4709 17911 4743
rect 18429 4573 18463 4607
rect 34069 4573 34103 4607
rect 18061 4505 18095 4539
rect 18613 4505 18647 4539
rect 1409 4437 1443 4471
rect 33701 4437 33735 4471
rect 34253 4437 34287 4471
rect 1409 4097 1443 4131
rect 1869 4097 1903 4131
rect 33425 4097 33459 4131
rect 34069 4097 34103 4131
rect 1593 3961 1627 3995
rect 2053 3893 2087 3927
rect 2329 3893 2363 3927
rect 33793 3893 33827 3927
rect 34253 3893 34287 3927
rect 8125 3689 8159 3723
rect 18337 3689 18371 3723
rect 32873 3689 32907 3723
rect 2145 3621 2179 3655
rect 2513 3621 2547 3655
rect 18061 3621 18095 3655
rect 33701 3621 33735 3655
rect 34069 3553 34103 3587
rect 1685 3485 1719 3519
rect 1961 3485 1995 3519
rect 2697 3485 2731 3519
rect 16681 3485 16715 3519
rect 17877 3485 17911 3519
rect 18521 3485 18555 3519
rect 32413 3485 32447 3519
rect 33505 3485 33539 3519
rect 19625 3417 19659 3451
rect 34253 3417 34287 3451
rect 1501 3349 1535 3383
rect 2973 3349 3007 3383
rect 3801 3349 3835 3383
rect 4169 3349 4203 3383
rect 16865 3349 16899 3383
rect 19349 3349 19383 3383
rect 33149 3349 33183 3383
rect 8033 3145 8067 3179
rect 13645 3145 13679 3179
rect 18981 3145 19015 3179
rect 22017 3145 22051 3179
rect 22845 3145 22879 3179
rect 25145 3145 25179 3179
rect 29745 3145 29779 3179
rect 17877 3077 17911 3111
rect 18705 3077 18739 3111
rect 1961 3009 1995 3043
rect 2513 3009 2547 3043
rect 4261 3009 4295 3043
rect 6837 3009 6871 3043
rect 7849 3009 7883 3043
rect 8677 3009 8711 3043
rect 11621 3009 11655 3043
rect 13829 3009 13863 3043
rect 14381 3009 14415 3043
rect 17141 3009 17175 3043
rect 17417 3009 17451 3043
rect 18061 3009 18095 3043
rect 18521 3009 18555 3043
rect 19165 3009 19199 3043
rect 19717 3009 19751 3043
rect 20177 3009 20211 3043
rect 22201 3009 22235 3043
rect 22477 3009 22511 3043
rect 24869 3009 24903 3043
rect 27445 3009 27479 3043
rect 27721 3009 27755 3043
rect 29929 3009 29963 3043
rect 30205 3009 30239 3043
rect 32321 3009 32355 3043
rect 32965 3009 32999 3043
rect 33793 3009 33827 3043
rect 2237 2941 2271 2975
rect 8309 2941 8343 2975
rect 31769 2941 31803 2975
rect 33517 2941 33551 2975
rect 3065 2873 3099 2907
rect 8861 2873 8895 2907
rect 12081 2873 12115 2907
rect 14197 2873 14231 2907
rect 17601 2873 17635 2907
rect 19993 2873 20027 2907
rect 31309 2873 31343 2907
rect 2697 2805 2731 2839
rect 3433 2805 3467 2839
rect 4077 2805 4111 2839
rect 4721 2805 4755 2839
rect 5917 2805 5951 2839
rect 6653 2805 6687 2839
rect 9137 2805 9171 2839
rect 11805 2805 11839 2839
rect 13369 2805 13403 2839
rect 14657 2805 14691 2839
rect 16957 2805 16991 2839
rect 19533 2805 19567 2839
rect 24685 2805 24719 2839
rect 27261 2805 27295 2839
rect 29469 2805 29503 2839
rect 32505 2805 32539 2839
rect 33149 2805 33183 2839
rect 14933 2601 14967 2635
rect 16313 2601 16347 2635
rect 23305 2601 23339 2635
rect 28641 2601 28675 2635
rect 31585 2533 31619 2567
rect 32965 2533 32999 2567
rect 2237 2465 2271 2499
rect 5181 2465 5215 2499
rect 6653 2465 6687 2499
rect 9413 2465 9447 2499
rect 18613 2465 18647 2499
rect 19257 2465 19291 2499
rect 19533 2465 19567 2499
rect 27261 2465 27295 2499
rect 29837 2465 29871 2499
rect 33517 2465 33551 2499
rect 1961 2397 1995 2431
rect 2789 2397 2823 2431
rect 3341 2397 3375 2431
rect 3801 2397 3835 2431
rect 4077 2397 4111 2431
rect 4905 2397 4939 2431
rect 6377 2397 6411 2431
rect 7757 2397 7791 2431
rect 8309 2397 8343 2431
rect 9137 2397 9171 2431
rect 10241 2397 10275 2431
rect 10977 2397 11011 2431
rect 11989 2397 12023 2431
rect 12633 2397 12667 2431
rect 13461 2397 13495 2431
rect 13737 2397 13771 2431
rect 14289 2397 14323 2431
rect 15117 2397 15151 2431
rect 15393 2397 15427 2431
rect 15853 2397 15887 2431
rect 16129 2397 16163 2431
rect 16957 2397 16991 2431
rect 17509 2397 17543 2431
rect 18889 2397 18923 2431
rect 20637 2397 20671 2431
rect 20913 2397 20947 2431
rect 22109 2397 22143 2431
rect 22937 2397 22971 2431
rect 23489 2397 23523 2431
rect 23765 2397 23799 2431
rect 24409 2397 24443 2431
rect 25237 2397 25271 2431
rect 26985 2397 27019 2431
rect 28089 2397 28123 2431
rect 28825 2397 28859 2431
rect 29561 2397 29595 2431
rect 30941 2397 30975 2431
rect 31309 2397 31343 2431
rect 31769 2397 31803 2431
rect 32413 2397 32447 2431
rect 33793 2397 33827 2431
rect 2605 2329 2639 2363
rect 29101 2329 29135 2363
rect 33149 2329 33183 2363
rect 3157 2261 3191 2295
rect 7573 2261 7607 2295
rect 8493 2261 8527 2295
rect 10425 2261 10459 2295
rect 11161 2261 11195 2295
rect 11805 2261 11839 2295
rect 12449 2261 12483 2295
rect 14473 2261 14507 2295
rect 16773 2261 16807 2295
rect 17693 2261 17727 2295
rect 20453 2261 20487 2295
rect 21925 2261 21959 2295
rect 22753 2261 22787 2295
rect 24593 2261 24627 2295
rect 25421 2261 25455 2295
rect 26525 2261 26559 2295
rect 28273 2261 28307 2295
rect 30757 2261 30791 2295
rect 32597 2261 32631 2295
<< metal1 >>
rect 11606 33940 11612 33992
rect 11664 33980 11670 33992
rect 18414 33980 18420 33992
rect 11664 33952 18420 33980
rect 11664 33940 11670 33952
rect 18414 33940 18420 33952
rect 18472 33940 18478 33992
rect 10502 33872 10508 33924
rect 10560 33912 10566 33924
rect 15010 33912 15016 33924
rect 10560 33884 15016 33912
rect 10560 33872 10566 33884
rect 15010 33872 15016 33884
rect 15068 33872 15074 33924
rect 16666 33872 16672 33924
rect 16724 33912 16730 33924
rect 20254 33912 20260 33924
rect 16724 33884 20260 33912
rect 16724 33872 16730 33884
rect 20254 33872 20260 33884
rect 20312 33872 20318 33924
rect 14366 33804 14372 33856
rect 14424 33844 14430 33856
rect 18966 33844 18972 33856
rect 14424 33816 18972 33844
rect 14424 33804 14430 33816
rect 18966 33804 18972 33816
rect 19024 33804 19030 33856
rect 1104 33754 34868 33776
rect 1104 33702 12214 33754
rect 12266 33702 12278 33754
rect 12330 33702 12342 33754
rect 12394 33702 12406 33754
rect 12458 33702 12470 33754
rect 12522 33702 23478 33754
rect 23530 33702 23542 33754
rect 23594 33702 23606 33754
rect 23658 33702 23670 33754
rect 23722 33702 23734 33754
rect 23786 33702 34868 33754
rect 1104 33680 34868 33702
rect 3878 33600 3884 33652
rect 3936 33640 3942 33652
rect 4157 33643 4215 33649
rect 4157 33640 4169 33643
rect 3936 33612 4169 33640
rect 3936 33600 3942 33612
rect 4157 33609 4169 33612
rect 4203 33609 4215 33643
rect 6730 33640 6736 33652
rect 6691 33612 6736 33640
rect 4157 33603 4215 33609
rect 6730 33600 6736 33612
rect 6788 33600 6794 33652
rect 9858 33640 9864 33652
rect 9819 33612 9864 33640
rect 9858 33600 9864 33612
rect 9916 33600 9922 33652
rect 16666 33640 16672 33652
rect 9968 33612 16672 33640
rect 2774 33572 2780 33584
rect 2735 33544 2780 33572
rect 2774 33532 2780 33544
rect 2832 33572 2838 33584
rect 3237 33575 3295 33581
rect 3237 33572 3249 33575
rect 2832 33544 3249 33572
rect 2832 33532 2838 33544
rect 3237 33541 3249 33544
rect 3283 33541 3295 33575
rect 9968 33572 9996 33612
rect 16666 33600 16672 33612
rect 16724 33600 16730 33652
rect 16758 33600 16764 33652
rect 16816 33640 16822 33652
rect 16945 33643 17003 33649
rect 16945 33640 16957 33643
rect 16816 33612 16957 33640
rect 16816 33600 16822 33612
rect 16945 33609 16957 33612
rect 16991 33609 17003 33643
rect 16945 33603 17003 33609
rect 18046 33600 18052 33652
rect 18104 33640 18110 33652
rect 18233 33643 18291 33649
rect 18233 33640 18245 33643
rect 18104 33612 18245 33640
rect 18104 33600 18110 33612
rect 18233 33609 18245 33612
rect 18279 33609 18291 33643
rect 23014 33640 23020 33652
rect 22975 33612 23020 33640
rect 18233 33603 18291 33609
rect 23014 33600 23020 33612
rect 23072 33600 23078 33652
rect 23934 33640 23940 33652
rect 23895 33612 23940 33640
rect 23934 33600 23940 33612
rect 23992 33600 23998 33652
rect 26050 33640 26056 33652
rect 26011 33612 26056 33640
rect 26050 33600 26056 33612
rect 26108 33600 26114 33652
rect 26510 33640 26516 33652
rect 26471 33612 26516 33640
rect 26510 33600 26516 33612
rect 26568 33600 26574 33652
rect 28166 33640 28172 33652
rect 28127 33612 28172 33640
rect 28166 33600 28172 33612
rect 28224 33600 28230 33652
rect 29086 33640 29092 33652
rect 29047 33612 29092 33640
rect 29086 33600 29092 33612
rect 29144 33600 29150 33652
rect 29914 33640 29920 33652
rect 29875 33612 29920 33640
rect 29914 33600 29920 33612
rect 29972 33600 29978 33652
rect 31754 33640 31760 33652
rect 31715 33612 31760 33640
rect 31754 33600 31760 33612
rect 31812 33600 31818 33652
rect 14734 33572 14740 33584
rect 3237 33535 3295 33541
rect 3896 33544 9996 33572
rect 10060 33544 14740 33572
rect 1026 33464 1032 33516
rect 1084 33504 1090 33516
rect 2222 33504 2228 33516
rect 1084 33476 2228 33504
rect 1084 33464 1090 33476
rect 2222 33464 2228 33476
rect 2280 33464 2286 33516
rect 2961 33507 3019 33513
rect 2961 33473 2973 33507
rect 3007 33504 3019 33507
rect 3896 33504 3924 33544
rect 3007 33476 3924 33504
rect 3007 33473 3019 33476
rect 2961 33467 3019 33473
rect 3970 33464 3976 33516
rect 4028 33504 4034 33516
rect 4614 33504 4620 33516
rect 4028 33476 4073 33504
rect 4575 33476 4620 33504
rect 4028 33464 4034 33476
rect 4614 33464 4620 33476
rect 4672 33464 4678 33516
rect 5534 33464 5540 33516
rect 5592 33504 5598 33516
rect 5721 33507 5779 33513
rect 5721 33504 5733 33507
rect 5592 33476 5733 33504
rect 5592 33464 5598 33476
rect 5721 33473 5733 33476
rect 5767 33473 5779 33507
rect 5721 33467 5779 33473
rect 6362 33464 6368 33516
rect 6420 33504 6426 33516
rect 6549 33507 6607 33513
rect 6549 33504 6561 33507
rect 6420 33476 6561 33504
rect 6420 33464 6426 33476
rect 6549 33473 6561 33476
rect 6595 33473 6607 33507
rect 7926 33504 7932 33516
rect 7887 33476 7932 33504
rect 6549 33467 6607 33473
rect 7926 33464 7932 33476
rect 7984 33504 7990 33516
rect 8389 33507 8447 33513
rect 8389 33504 8401 33507
rect 7984 33476 8401 33504
rect 7984 33464 7990 33476
rect 8389 33473 8401 33476
rect 8435 33473 8447 33507
rect 8389 33467 8447 33473
rect 8478 33464 8484 33516
rect 8536 33504 8542 33516
rect 10060 33513 10088 33544
rect 14734 33532 14740 33544
rect 14792 33532 14798 33584
rect 15470 33532 15476 33584
rect 15528 33572 15534 33584
rect 17405 33575 17463 33581
rect 17405 33572 17417 33575
rect 15528 33544 17417 33572
rect 15528 33532 15534 33544
rect 9217 33507 9275 33513
rect 9217 33504 9229 33507
rect 8536 33476 9229 33504
rect 8536 33464 8542 33476
rect 9217 33473 9229 33476
rect 9263 33473 9275 33507
rect 9217 33467 9275 33473
rect 10045 33507 10103 33513
rect 10045 33473 10057 33507
rect 10091 33473 10103 33507
rect 10045 33467 10103 33473
rect 10873 33507 10931 33513
rect 10873 33473 10885 33507
rect 10919 33504 10931 33507
rect 11698 33504 11704 33516
rect 10919 33476 11560 33504
rect 11659 33476 11704 33504
rect 10919 33473 10931 33476
rect 10873 33467 10931 33473
rect 1949 33439 2007 33445
rect 1949 33405 1961 33439
rect 1995 33405 2007 33439
rect 1949 33399 2007 33405
rect 1964 33368 1992 33399
rect 3050 33396 3056 33448
rect 3108 33436 3114 33448
rect 4893 33439 4951 33445
rect 4893 33436 4905 33439
rect 3108 33408 4905 33436
rect 3108 33396 3114 33408
rect 4893 33405 4905 33408
rect 4939 33405 4951 33439
rect 10502 33436 10508 33448
rect 4893 33399 4951 33405
rect 5000 33408 10508 33436
rect 5000 33368 5028 33408
rect 10502 33396 10508 33408
rect 10560 33396 10566 33448
rect 10594 33396 10600 33448
rect 10652 33436 10658 33448
rect 11146 33436 11152 33448
rect 10652 33408 11152 33436
rect 10652 33396 10658 33408
rect 11146 33396 11152 33408
rect 11204 33396 11210 33448
rect 11532 33436 11560 33476
rect 11698 33464 11704 33476
rect 11756 33504 11762 33516
rect 12161 33507 12219 33513
rect 12161 33504 12173 33507
rect 11756 33476 12173 33504
rect 11756 33464 11762 33476
rect 12161 33473 12173 33476
rect 12207 33473 12219 33507
rect 12161 33467 12219 33473
rect 13725 33507 13783 33513
rect 13725 33473 13737 33507
rect 13771 33504 13783 33507
rect 14366 33504 14372 33516
rect 13771 33476 14372 33504
rect 13771 33473 13783 33476
rect 13725 33467 13783 33473
rect 14366 33464 14372 33476
rect 14424 33464 14430 33516
rect 14458 33464 14464 33516
rect 14516 33504 14522 33516
rect 14645 33507 14703 33513
rect 14645 33504 14657 33507
rect 14516 33476 14657 33504
rect 14516 33464 14522 33476
rect 14645 33473 14657 33476
rect 14691 33504 14703 33507
rect 15105 33507 15163 33513
rect 15105 33504 15117 33507
rect 14691 33476 15117 33504
rect 14691 33473 14703 33476
rect 14645 33467 14703 33473
rect 15105 33473 15117 33476
rect 15151 33473 15163 33507
rect 15105 33467 15163 33473
rect 15948 33436 15976 33544
rect 17405 33541 17417 33544
rect 17451 33541 17463 33575
rect 17405 33535 17463 33541
rect 18598 33532 18604 33584
rect 18656 33572 18662 33584
rect 18656 33544 20944 33572
rect 18656 33532 18662 33544
rect 16025 33507 16083 33513
rect 16025 33473 16037 33507
rect 16071 33504 16083 33507
rect 17126 33504 17132 33516
rect 16071 33476 16574 33504
rect 17087 33476 17132 33504
rect 16071 33473 16083 33476
rect 16025 33467 16083 33473
rect 16301 33439 16359 33445
rect 16301 33436 16313 33439
rect 11532 33408 15792 33436
rect 15948 33408 16313 33436
rect 1964 33340 5028 33368
rect 5905 33371 5963 33377
rect 5905 33337 5917 33371
rect 5951 33368 5963 33371
rect 11606 33368 11612 33380
rect 5951 33340 11612 33368
rect 5951 33337 5963 33340
rect 5905 33331 5963 33337
rect 11606 33328 11612 33340
rect 11664 33328 11670 33380
rect 11716 33340 13768 33368
rect 2590 33260 2596 33312
rect 2648 33300 2654 33312
rect 3970 33300 3976 33312
rect 2648 33272 3976 33300
rect 2648 33260 2654 33272
rect 3970 33260 3976 33272
rect 4028 33260 4034 33312
rect 8018 33300 8024 33312
rect 7979 33272 8024 33300
rect 8018 33260 8024 33272
rect 8076 33260 8082 33312
rect 9309 33303 9367 33309
rect 9309 33269 9321 33303
rect 9355 33300 9367 33303
rect 11716 33300 11744 33340
rect 11882 33300 11888 33312
rect 9355 33272 11744 33300
rect 11843 33272 11888 33300
rect 9355 33269 9367 33272
rect 9309 33263 9367 33269
rect 11882 33260 11888 33272
rect 11940 33260 11946 33312
rect 13740 33300 13768 33340
rect 13814 33328 13820 33380
rect 13872 33368 13878 33380
rect 14185 33371 14243 33377
rect 14185 33368 14197 33371
rect 13872 33340 14197 33368
rect 13872 33328 13878 33340
rect 14185 33337 14197 33340
rect 14231 33337 14243 33371
rect 14185 33331 14243 33337
rect 14829 33371 14887 33377
rect 14829 33337 14841 33371
rect 14875 33368 14887 33371
rect 15764 33368 15792 33408
rect 16301 33405 16313 33408
rect 16347 33405 16359 33439
rect 16546 33436 16574 33476
rect 17126 33464 17132 33476
rect 17184 33464 17190 33516
rect 18417 33507 18475 33513
rect 18417 33473 18429 33507
rect 18463 33504 18475 33507
rect 18782 33504 18788 33516
rect 18463 33476 18788 33504
rect 18463 33473 18475 33476
rect 18417 33467 18475 33473
rect 18782 33464 18788 33476
rect 18840 33464 18846 33516
rect 18877 33507 18935 33513
rect 18877 33473 18889 33507
rect 18923 33504 18935 33507
rect 19426 33504 19432 33516
rect 18923 33476 19432 33504
rect 18923 33473 18935 33476
rect 18877 33467 18935 33473
rect 19426 33464 19432 33476
rect 19484 33464 19490 33516
rect 20622 33504 20628 33516
rect 20583 33476 20628 33504
rect 20622 33464 20628 33476
rect 20680 33464 20686 33516
rect 20916 33513 20944 33544
rect 20901 33507 20959 33513
rect 20901 33473 20913 33507
rect 20947 33473 20959 33507
rect 20901 33467 20959 33473
rect 21266 33464 21272 33516
rect 21324 33504 21330 33516
rect 21821 33507 21879 33513
rect 21821 33504 21833 33507
rect 21324 33476 21833 33504
rect 21324 33464 21330 33476
rect 21821 33473 21833 33476
rect 21867 33504 21879 33507
rect 22281 33507 22339 33513
rect 22281 33504 22293 33507
rect 21867 33476 22293 33504
rect 21867 33473 21879 33476
rect 21821 33467 21879 33473
rect 22281 33473 22293 33476
rect 22327 33473 22339 33507
rect 23032 33504 23060 33600
rect 23477 33507 23535 33513
rect 23477 33504 23489 33507
rect 23032 33476 23489 33504
rect 22281 33467 22339 33473
rect 23477 33473 23489 33476
rect 23523 33473 23535 33507
rect 23952 33504 23980 33600
rect 24397 33507 24455 33513
rect 24397 33504 24409 33507
rect 23952 33476 24409 33504
rect 23477 33467 23535 33473
rect 24397 33473 24409 33476
rect 24443 33473 24455 33507
rect 24397 33467 24455 33473
rect 25593 33507 25651 33513
rect 25593 33473 25605 33507
rect 25639 33504 25651 33507
rect 25866 33504 25872 33516
rect 25639 33476 25872 33504
rect 25639 33473 25651 33476
rect 25593 33467 25651 33473
rect 25866 33464 25872 33476
rect 25924 33464 25930 33516
rect 26528 33504 26556 33600
rect 26973 33507 27031 33513
rect 26973 33504 26985 33507
rect 26528 33476 26985 33504
rect 26973 33473 26985 33476
rect 27019 33473 27031 33507
rect 28184 33504 28212 33600
rect 31772 33572 31800 33600
rect 32493 33575 32551 33581
rect 32493 33572 32505 33575
rect 31772 33544 32505 33572
rect 32493 33541 32505 33544
rect 32539 33541 32551 33575
rect 32493 33535 32551 33541
rect 28445 33507 28503 33513
rect 28445 33504 28457 33507
rect 28184 33476 28457 33504
rect 26973 33467 27031 33473
rect 28445 33473 28457 33476
rect 28491 33473 28503 33507
rect 28445 33467 28503 33473
rect 28718 33464 28724 33516
rect 28776 33504 28782 33516
rect 28905 33507 28963 33513
rect 28905 33504 28917 33507
rect 28776 33476 28917 33504
rect 28776 33464 28782 33476
rect 28905 33473 28917 33476
rect 28951 33473 28963 33507
rect 28905 33467 28963 33473
rect 29733 33507 29791 33513
rect 29733 33473 29745 33507
rect 29779 33473 29791 33507
rect 30374 33504 30380 33516
rect 30335 33476 30380 33504
rect 29733 33467 29791 33473
rect 17402 33436 17408 33448
rect 16546 33408 17408 33436
rect 16301 33399 16359 33405
rect 17402 33396 17408 33408
rect 17460 33396 17466 33448
rect 19705 33439 19763 33445
rect 19705 33405 19717 33439
rect 19751 33436 19763 33439
rect 19794 33436 19800 33448
rect 19751 33408 19800 33436
rect 19751 33405 19763 33408
rect 19705 33399 19763 33405
rect 19794 33396 19800 33408
rect 19852 33396 19858 33448
rect 24486 33396 24492 33448
rect 24544 33436 24550 33448
rect 24673 33439 24731 33445
rect 24673 33436 24685 33439
rect 24544 33408 24685 33436
rect 24544 33396 24550 33408
rect 24673 33405 24685 33408
rect 24719 33405 24731 33439
rect 24673 33399 24731 33405
rect 27249 33439 27307 33445
rect 27249 33405 27261 33439
rect 27295 33436 27307 33439
rect 27338 33436 27344 33448
rect 27295 33408 27344 33436
rect 27295 33405 27307 33408
rect 27249 33399 27307 33405
rect 27338 33396 27344 33408
rect 27396 33396 27402 33448
rect 27614 33396 27620 33448
rect 27672 33436 27678 33448
rect 29748 33436 29776 33467
rect 30374 33464 30380 33476
rect 30432 33464 30438 33516
rect 33137 33507 33195 33513
rect 33137 33473 33149 33507
rect 33183 33504 33195 33507
rect 33318 33504 33324 33516
rect 33183 33476 33324 33504
rect 33183 33473 33195 33476
rect 33137 33467 33195 33473
rect 33318 33464 33324 33476
rect 33376 33504 33382 33516
rect 34422 33504 34428 33516
rect 33376 33476 34428 33504
rect 33376 33464 33382 33476
rect 34422 33464 34428 33476
rect 34480 33464 34486 33516
rect 27672 33408 29776 33436
rect 30653 33439 30711 33445
rect 27672 33396 27678 33408
rect 30653 33405 30665 33439
rect 30699 33436 30711 33439
rect 31202 33436 31208 33448
rect 30699 33408 31208 33436
rect 30699 33405 30711 33408
rect 30653 33399 30711 33405
rect 31202 33396 31208 33408
rect 31260 33396 31266 33448
rect 33226 33396 33232 33448
rect 33284 33436 33290 33448
rect 33505 33439 33563 33445
rect 33505 33436 33517 33439
rect 33284 33408 33517 33436
rect 33284 33396 33290 33408
rect 33505 33405 33517 33408
rect 33551 33436 33563 33439
rect 33594 33436 33600 33448
rect 33551 33408 33600 33436
rect 33551 33405 33563 33408
rect 33505 33399 33563 33405
rect 33594 33396 33600 33408
rect 33652 33396 33658 33448
rect 33778 33436 33784 33448
rect 33739 33408 33784 33436
rect 33778 33396 33784 33408
rect 33836 33396 33842 33448
rect 17770 33368 17776 33380
rect 14875 33340 15700 33368
rect 15764 33340 17776 33368
rect 14875 33337 14887 33340
rect 14829 33331 14887 33337
rect 15562 33300 15568 33312
rect 13740 33272 15568 33300
rect 15562 33260 15568 33272
rect 15620 33260 15626 33312
rect 15672 33300 15700 33340
rect 17770 33328 17776 33340
rect 17828 33328 17834 33380
rect 19334 33328 19340 33380
rect 19392 33368 19398 33380
rect 23293 33371 23351 33377
rect 23293 33368 23305 33371
rect 19392 33340 23305 33368
rect 19392 33328 19398 33340
rect 23293 33337 23305 33340
rect 23339 33337 23351 33371
rect 32306 33368 32312 33380
rect 32267 33340 32312 33368
rect 23293 33331 23351 33337
rect 32306 33328 32312 33340
rect 32364 33328 32370 33380
rect 32858 33328 32864 33380
rect 32916 33368 32922 33380
rect 32953 33371 33011 33377
rect 32953 33368 32965 33371
rect 32916 33340 32965 33368
rect 32916 33328 32922 33340
rect 32953 33337 32965 33340
rect 32999 33337 33011 33371
rect 32953 33331 33011 33337
rect 18506 33300 18512 33312
rect 15672 33272 18512 33300
rect 18506 33260 18512 33272
rect 18564 33260 18570 33312
rect 21910 33260 21916 33312
rect 21968 33300 21974 33312
rect 22005 33303 22063 33309
rect 22005 33300 22017 33303
rect 21968 33272 22017 33300
rect 21968 33260 21974 33272
rect 22005 33269 22017 33272
rect 22051 33269 22063 33303
rect 22005 33263 22063 33269
rect 28629 33303 28687 33309
rect 28629 33269 28641 33303
rect 28675 33300 28687 33303
rect 30834 33300 30840 33312
rect 28675 33272 30840 33300
rect 28675 33269 28687 33272
rect 28629 33263 28687 33269
rect 30834 33260 30840 33272
rect 30892 33260 30898 33312
rect 1104 33210 34868 33232
rect 1104 33158 6582 33210
rect 6634 33158 6646 33210
rect 6698 33158 6710 33210
rect 6762 33158 6774 33210
rect 6826 33158 6838 33210
rect 6890 33158 17846 33210
rect 17898 33158 17910 33210
rect 17962 33158 17974 33210
rect 18026 33158 18038 33210
rect 18090 33158 18102 33210
rect 18154 33158 29110 33210
rect 29162 33158 29174 33210
rect 29226 33158 29238 33210
rect 29290 33158 29302 33210
rect 29354 33158 29366 33210
rect 29418 33158 34868 33210
rect 1104 33136 34868 33158
rect 2222 33056 2228 33108
rect 2280 33096 2286 33108
rect 2777 33099 2835 33105
rect 2777 33096 2789 33099
rect 2280 33068 2789 33096
rect 2280 33056 2286 33068
rect 2777 33065 2789 33068
rect 2823 33065 2835 33099
rect 2777 33059 2835 33065
rect 4525 33099 4583 33105
rect 4525 33065 4537 33099
rect 4571 33096 4583 33099
rect 4614 33096 4620 33108
rect 4571 33068 4620 33096
rect 4571 33065 4583 33068
rect 4525 33059 4583 33065
rect 4614 33056 4620 33068
rect 4672 33056 4678 33108
rect 5534 33096 5540 33108
rect 5495 33068 5540 33096
rect 5534 33056 5540 33068
rect 5592 33056 5598 33108
rect 5994 33096 6000 33108
rect 5955 33068 6000 33096
rect 5994 33056 6000 33068
rect 6052 33056 6058 33108
rect 8478 33096 8484 33108
rect 8439 33068 8484 33096
rect 8478 33056 8484 33068
rect 8536 33056 8542 33108
rect 10778 33096 10784 33108
rect 10739 33068 10784 33096
rect 10778 33056 10784 33068
rect 10836 33056 10842 33108
rect 11146 33056 11152 33108
rect 11204 33096 11210 33108
rect 11517 33099 11575 33105
rect 11517 33096 11529 33099
rect 11204 33068 11529 33096
rect 11204 33056 11210 33068
rect 11517 33065 11529 33068
rect 11563 33065 11575 33099
rect 14642 33096 14648 33108
rect 14603 33068 14648 33096
rect 11517 33059 11575 33065
rect 14642 33056 14648 33068
rect 14700 33056 14706 33108
rect 16390 33096 16396 33108
rect 16351 33068 16396 33096
rect 16390 33056 16396 33068
rect 16448 33056 16454 33108
rect 16945 33099 17003 33105
rect 16945 33065 16957 33099
rect 16991 33096 17003 33099
rect 17126 33096 17132 33108
rect 16991 33068 17132 33096
rect 16991 33065 17003 33068
rect 16945 33059 17003 33065
rect 17126 33056 17132 33068
rect 17184 33056 17190 33108
rect 18690 33056 18696 33108
rect 18748 33096 18754 33108
rect 19429 33099 19487 33105
rect 19429 33096 19441 33099
rect 18748 33068 19441 33096
rect 18748 33056 18754 33068
rect 19429 33065 19441 33068
rect 19475 33065 19487 33099
rect 19429 33059 19487 33065
rect 20622 33056 20628 33108
rect 20680 33096 20686 33108
rect 21545 33099 21603 33105
rect 21545 33096 21557 33099
rect 20680 33068 21557 33096
rect 20680 33056 20686 33068
rect 21545 33065 21557 33068
rect 21591 33065 21603 33099
rect 24670 33096 24676 33108
rect 21545 33059 21603 33065
rect 22020 33068 24532 33096
rect 24631 33068 24676 33096
rect 1302 32988 1308 33040
rect 1360 33028 1366 33040
rect 3145 33031 3203 33037
rect 3145 33028 3157 33031
rect 1360 33000 3157 33028
rect 1360 32988 1366 33000
rect 3145 32997 3157 33000
rect 3191 32997 3203 33031
rect 3145 32991 3203 32997
rect 14660 32960 14688 33056
rect 14734 32988 14740 33040
rect 14792 33028 14798 33040
rect 17405 33031 17463 33037
rect 17405 33028 17417 33031
rect 14792 33000 17417 33028
rect 14792 32988 14798 33000
rect 17405 32997 17417 33000
rect 17451 32997 17463 33031
rect 22020 33028 22048 33068
rect 17405 32991 17463 32997
rect 17604 33000 22048 33028
rect 22097 33031 22155 33037
rect 14921 32963 14979 32969
rect 14921 32960 14933 32963
rect 14660 32932 14933 32960
rect 14921 32929 14933 32932
rect 14967 32929 14979 32963
rect 14921 32923 14979 32929
rect 15010 32920 15016 32972
rect 15068 32960 15074 32972
rect 15068 32932 16574 32960
rect 15068 32920 15074 32932
rect 14 32852 20 32904
rect 72 32892 78 32904
rect 1302 32892 1308 32904
rect 72 32864 1308 32892
rect 72 32852 78 32864
rect 1302 32852 1308 32864
rect 1360 32892 1366 32904
rect 1673 32895 1731 32901
rect 1673 32892 1685 32895
rect 1360 32864 1685 32892
rect 1360 32852 1366 32864
rect 1673 32861 1685 32864
rect 1719 32861 1731 32895
rect 1673 32855 1731 32861
rect 2130 32852 2136 32904
rect 2188 32892 2194 32904
rect 2225 32895 2283 32901
rect 2225 32892 2237 32895
rect 2188 32864 2237 32892
rect 2188 32852 2194 32864
rect 2225 32861 2237 32864
rect 2271 32892 2283 32895
rect 2774 32892 2780 32904
rect 2271 32864 2780 32892
rect 2271 32861 2283 32864
rect 2225 32855 2283 32861
rect 2774 32852 2780 32864
rect 2832 32852 2838 32904
rect 3329 32895 3387 32901
rect 3329 32861 3341 32895
rect 3375 32892 3387 32895
rect 3510 32892 3516 32904
rect 3375 32864 3516 32892
rect 3375 32861 3387 32864
rect 3329 32855 3387 32861
rect 3510 32852 3516 32864
rect 3568 32852 3574 32904
rect 6181 32895 6239 32901
rect 6181 32861 6193 32895
rect 6227 32892 6239 32895
rect 9306 32892 9312 32904
rect 6227 32864 6500 32892
rect 9267 32864 9312 32892
rect 6227 32861 6239 32864
rect 6181 32855 6239 32861
rect 1854 32824 1860 32836
rect 1815 32796 1860 32824
rect 1854 32784 1860 32796
rect 1912 32784 1918 32836
rect 6472 32768 6500 32864
rect 9306 32852 9312 32864
rect 9364 32892 9370 32904
rect 9585 32895 9643 32901
rect 9585 32892 9597 32895
rect 9364 32864 9597 32892
rect 9364 32852 9370 32864
rect 9585 32861 9597 32864
rect 9631 32861 9643 32895
rect 9585 32855 9643 32861
rect 10778 32852 10784 32904
rect 10836 32892 10842 32904
rect 11057 32895 11115 32901
rect 11057 32892 11069 32895
rect 10836 32864 11069 32892
rect 10836 32852 10842 32864
rect 11057 32861 11069 32864
rect 11103 32861 11115 32895
rect 15194 32892 15200 32904
rect 15155 32864 15200 32892
rect 11057 32855 11115 32861
rect 15194 32852 15200 32864
rect 15252 32852 15258 32904
rect 15562 32852 15568 32904
rect 15620 32892 15626 32904
rect 16209 32895 16267 32901
rect 16209 32892 16221 32895
rect 15620 32864 16221 32892
rect 15620 32852 15626 32864
rect 16209 32861 16221 32864
rect 16255 32861 16267 32895
rect 16546 32892 16574 32932
rect 17604 32901 17632 33000
rect 22097 32997 22109 33031
rect 22143 32997 22155 33031
rect 24504 33028 24532 33068
rect 24670 33056 24676 33068
rect 24728 33056 24734 33108
rect 25406 33096 25412 33108
rect 25367 33068 25412 33096
rect 25406 33056 25412 33068
rect 25464 33056 25470 33108
rect 27246 33096 27252 33108
rect 27207 33068 27252 33096
rect 27246 33056 27252 33068
rect 27304 33056 27310 33108
rect 30285 33099 30343 33105
rect 27356 33068 27844 33096
rect 27356 33028 27384 33068
rect 24504 33000 27384 33028
rect 27709 33031 27767 33037
rect 22097 32991 22155 32997
rect 27709 32997 27721 33031
rect 27755 32997 27767 33031
rect 27816 33028 27844 33068
rect 30285 33065 30297 33099
rect 30331 33096 30343 33099
rect 30374 33096 30380 33108
rect 30331 33068 30380 33096
rect 30331 33065 30343 33068
rect 30285 33059 30343 33065
rect 30374 33056 30380 33068
rect 30432 33056 30438 33108
rect 30742 33096 30748 33108
rect 30703 33068 30748 33096
rect 30742 33056 30748 33068
rect 30800 33056 30806 33108
rect 32490 33096 32496 33108
rect 32451 33068 32496 33096
rect 32490 33056 32496 33068
rect 32548 33056 32554 33108
rect 33134 33096 33140 33108
rect 33095 33068 33140 33096
rect 33134 33056 33140 33068
rect 33192 33056 33198 33108
rect 33686 33096 33692 33108
rect 33647 33068 33692 33096
rect 33686 33056 33692 33068
rect 33744 33056 33750 33108
rect 33778 33028 33784 33040
rect 27816 33000 33784 33028
rect 27709 32991 27767 32997
rect 16761 32895 16819 32901
rect 16761 32892 16773 32895
rect 16546 32864 16773 32892
rect 16209 32855 16267 32861
rect 16761 32861 16773 32864
rect 16807 32861 16819 32895
rect 16761 32855 16819 32861
rect 17589 32895 17647 32901
rect 17589 32861 17601 32895
rect 17635 32861 17647 32895
rect 17589 32855 17647 32861
rect 18049 32895 18107 32901
rect 18049 32861 18061 32895
rect 18095 32892 18107 32895
rect 19242 32892 19248 32904
rect 18095 32864 19104 32892
rect 19203 32864 19248 32892
rect 18095 32861 18107 32864
rect 18049 32855 18107 32861
rect 15286 32784 15292 32836
rect 15344 32824 15350 32836
rect 17865 32827 17923 32833
rect 17865 32824 17877 32827
rect 15344 32796 17877 32824
rect 15344 32784 15350 32796
rect 17865 32793 17877 32796
rect 17911 32793 17923 32827
rect 18506 32824 18512 32836
rect 18467 32796 18512 32824
rect 17865 32787 17923 32793
rect 18506 32784 18512 32796
rect 18564 32784 18570 32836
rect 19076 32824 19104 32864
rect 19242 32852 19248 32864
rect 19300 32852 19306 32904
rect 21910 32892 21916 32904
rect 21871 32864 21916 32892
rect 21910 32852 21916 32864
rect 21968 32852 21974 32904
rect 22112 32892 22140 32991
rect 27724 32960 27752 32991
rect 33778 32988 33784 33000
rect 33836 32988 33842 33040
rect 29914 32960 29920 32972
rect 24872 32932 27752 32960
rect 27816 32932 29920 32960
rect 24872 32901 24900 32932
rect 24857 32895 24915 32901
rect 22112 32864 24808 32892
rect 19334 32824 19340 32836
rect 19076 32796 19340 32824
rect 19334 32784 19340 32796
rect 19392 32784 19398 32836
rect 24780 32824 24808 32864
rect 24857 32861 24869 32895
rect 24903 32861 24915 32895
rect 24857 32855 24915 32861
rect 25225 32895 25283 32901
rect 25225 32861 25237 32895
rect 25271 32861 25283 32895
rect 25225 32855 25283 32861
rect 27433 32895 27491 32901
rect 27433 32861 27445 32895
rect 27479 32892 27491 32895
rect 27816 32892 27844 32932
rect 29914 32920 29920 32932
rect 29972 32920 29978 32972
rect 30742 32920 30748 32972
rect 30800 32960 30806 32972
rect 31021 32963 31079 32969
rect 31021 32960 31033 32963
rect 30800 32932 31033 32960
rect 30800 32920 30806 32932
rect 31021 32929 31033 32932
rect 31067 32929 31079 32963
rect 31021 32923 31079 32929
rect 31938 32920 31944 32972
rect 31996 32960 32002 32972
rect 31996 32932 33548 32960
rect 31996 32920 32002 32932
rect 27479 32888 27660 32892
rect 27724 32888 27844 32892
rect 27479 32864 27844 32888
rect 27479 32861 27491 32864
rect 27433 32855 27491 32861
rect 27632 32860 27752 32864
rect 25240 32824 25268 32855
rect 27890 32852 27896 32904
rect 27948 32892 27954 32904
rect 31294 32892 31300 32904
rect 27948 32864 27993 32892
rect 31255 32864 31300 32892
rect 27948 32852 27954 32864
rect 31294 32852 31300 32864
rect 31352 32852 31358 32904
rect 32309 32895 32367 32901
rect 32309 32861 32321 32895
rect 32355 32861 32367 32895
rect 32950 32892 32956 32904
rect 32911 32864 32956 32892
rect 32309 32855 32367 32861
rect 32324 32824 32352 32855
rect 32950 32852 32956 32864
rect 33008 32852 33014 32904
rect 33520 32901 33548 32932
rect 33505 32895 33563 32901
rect 33505 32861 33517 32895
rect 33551 32861 33563 32895
rect 34238 32892 34244 32904
rect 34199 32864 34244 32892
rect 33505 32855 33563 32861
rect 34238 32852 34244 32864
rect 34296 32852 34302 32904
rect 24780 32796 25268 32824
rect 28184 32796 32352 32824
rect 2314 32756 2320 32768
rect 2275 32728 2320 32756
rect 2314 32716 2320 32728
rect 2372 32716 2378 32768
rect 6454 32756 6460 32768
rect 6415 32728 6460 32756
rect 6454 32716 6460 32728
rect 6512 32716 6518 32768
rect 9122 32756 9128 32768
rect 9083 32728 9128 32756
rect 9122 32716 9128 32728
rect 9180 32716 9186 32768
rect 11238 32756 11244 32768
rect 11199 32728 11244 32756
rect 11238 32716 11244 32728
rect 11296 32716 11302 32768
rect 18601 32759 18659 32765
rect 18601 32725 18613 32759
rect 18647 32756 18659 32759
rect 28184 32756 28212 32796
rect 32766 32784 32772 32836
rect 32824 32824 32830 32836
rect 34256 32824 34284 32852
rect 32824 32796 34284 32824
rect 32824 32784 32830 32796
rect 28718 32756 28724 32768
rect 18647 32728 28212 32756
rect 28679 32728 28724 32756
rect 18647 32725 18659 32728
rect 18601 32719 18659 32725
rect 28718 32716 28724 32728
rect 28776 32716 28782 32768
rect 28810 32716 28816 32768
rect 28868 32756 28874 32768
rect 34149 32759 34207 32765
rect 34149 32756 34161 32759
rect 28868 32728 34161 32756
rect 28868 32716 28874 32728
rect 34149 32725 34161 32728
rect 34195 32725 34207 32759
rect 34149 32719 34207 32725
rect 1104 32666 34868 32688
rect 1104 32614 12214 32666
rect 12266 32614 12278 32666
rect 12330 32614 12342 32666
rect 12394 32614 12406 32666
rect 12458 32614 12470 32666
rect 12522 32614 23478 32666
rect 23530 32614 23542 32666
rect 23594 32614 23606 32666
rect 23658 32614 23670 32666
rect 23722 32614 23734 32666
rect 23786 32614 34868 32666
rect 1104 32592 34868 32614
rect 2593 32555 2651 32561
rect 2593 32521 2605 32555
rect 2639 32552 2651 32555
rect 2866 32552 2872 32564
rect 2639 32524 2872 32552
rect 2639 32521 2651 32524
rect 2593 32515 2651 32521
rect 2866 32512 2872 32524
rect 2924 32512 2930 32564
rect 15562 32552 15568 32564
rect 15523 32524 15568 32552
rect 15562 32512 15568 32524
rect 15620 32512 15626 32564
rect 24854 32512 24860 32564
rect 24912 32552 24918 32564
rect 28810 32552 28816 32564
rect 24912 32524 28816 32552
rect 24912 32512 24918 32524
rect 28810 32512 28816 32524
rect 28868 32512 28874 32564
rect 32766 32552 32772 32564
rect 32727 32524 32772 32552
rect 32766 32512 32772 32524
rect 32824 32512 32830 32564
rect 33045 32555 33103 32561
rect 33045 32521 33057 32555
rect 33091 32521 33103 32555
rect 33045 32515 33103 32521
rect 33689 32555 33747 32561
rect 33689 32521 33701 32555
rect 33735 32552 33747 32555
rect 34146 32552 34152 32564
rect 33735 32524 34152 32552
rect 33735 32521 33747 32524
rect 33689 32515 33747 32521
rect 1302 32444 1308 32496
rect 1360 32484 1366 32496
rect 3053 32487 3111 32493
rect 3053 32484 3065 32487
rect 1360 32456 3065 32484
rect 1360 32444 1366 32456
rect 3053 32453 3065 32456
rect 3099 32453 3111 32487
rect 17865 32487 17923 32493
rect 17865 32484 17877 32487
rect 3053 32447 3111 32453
rect 6886 32456 17877 32484
rect 2777 32419 2835 32425
rect 2777 32385 2789 32419
rect 2823 32416 2835 32419
rect 6886 32416 6914 32456
rect 17865 32453 17877 32456
rect 17911 32453 17923 32487
rect 17865 32447 17923 32453
rect 18049 32487 18107 32493
rect 18049 32453 18061 32487
rect 18095 32484 18107 32487
rect 18095 32456 22094 32484
rect 18095 32453 18107 32456
rect 18049 32447 18107 32453
rect 2823 32388 6914 32416
rect 2823 32385 2835 32388
rect 2777 32379 2835 32385
rect 11238 32376 11244 32428
rect 11296 32416 11302 32428
rect 15381 32419 15439 32425
rect 15381 32416 15393 32419
rect 11296 32388 15393 32416
rect 11296 32376 11302 32388
rect 15381 32385 15393 32388
rect 15427 32385 15439 32419
rect 18506 32416 18512 32428
rect 18467 32388 18512 32416
rect 15381 32379 15439 32385
rect 18506 32376 18512 32388
rect 18564 32416 18570 32428
rect 18969 32419 19027 32425
rect 18969 32416 18981 32419
rect 18564 32388 18981 32416
rect 18564 32376 18570 32388
rect 18969 32385 18981 32388
rect 19015 32385 19027 32419
rect 22066 32416 22094 32456
rect 27890 32444 27896 32496
rect 27948 32484 27954 32496
rect 33060 32484 33088 32515
rect 34146 32512 34152 32524
rect 34204 32512 34210 32564
rect 27948 32456 33088 32484
rect 27948 32444 27954 32456
rect 30374 32416 30380 32428
rect 22066 32388 30380 32416
rect 18969 32379 19027 32385
rect 30374 32376 30380 32388
rect 30432 32376 30438 32428
rect 33229 32419 33287 32425
rect 33229 32385 33241 32419
rect 33275 32416 33287 32419
rect 33410 32416 33416 32428
rect 33275 32388 33416 32416
rect 33275 32385 33287 32388
rect 33229 32379 33287 32385
rect 33410 32376 33416 32388
rect 33468 32376 33474 32428
rect 33505 32419 33563 32425
rect 33505 32385 33517 32419
rect 33551 32385 33563 32419
rect 33505 32379 33563 32385
rect 1394 32348 1400 32360
rect 1355 32320 1400 32348
rect 1394 32308 1400 32320
rect 1452 32308 1458 32360
rect 1673 32351 1731 32357
rect 1673 32317 1685 32351
rect 1719 32348 1731 32351
rect 1762 32348 1768 32360
rect 1719 32320 1768 32348
rect 1719 32317 1731 32320
rect 1673 32311 1731 32317
rect 1762 32308 1768 32320
rect 1820 32308 1826 32360
rect 32401 32351 32459 32357
rect 32401 32317 32413 32351
rect 32447 32348 32459 32351
rect 33318 32348 33324 32360
rect 32447 32320 33324 32348
rect 32447 32317 32459 32320
rect 32401 32311 32459 32317
rect 33318 32308 33324 32320
rect 33376 32308 33382 32360
rect 18693 32283 18751 32289
rect 18693 32249 18705 32283
rect 18739 32280 18751 32283
rect 33520 32280 33548 32379
rect 33594 32376 33600 32428
rect 33652 32416 33658 32428
rect 34057 32419 34115 32425
rect 34057 32416 34069 32419
rect 33652 32388 34069 32416
rect 33652 32376 33658 32388
rect 34057 32385 34069 32388
rect 34103 32385 34115 32419
rect 34057 32379 34115 32385
rect 18739 32252 33548 32280
rect 18739 32249 18751 32252
rect 18693 32243 18751 32249
rect 31757 32215 31815 32221
rect 31757 32181 31769 32215
rect 31803 32212 31815 32215
rect 31938 32212 31944 32224
rect 31803 32184 31944 32212
rect 31803 32181 31815 32184
rect 31757 32175 31815 32181
rect 31938 32172 31944 32184
rect 31996 32172 32002 32224
rect 34238 32212 34244 32224
rect 34199 32184 34244 32212
rect 34238 32172 34244 32184
rect 34296 32172 34302 32224
rect 1104 32122 34868 32144
rect 1104 32070 6582 32122
rect 6634 32070 6646 32122
rect 6698 32070 6710 32122
rect 6762 32070 6774 32122
rect 6826 32070 6838 32122
rect 6890 32070 17846 32122
rect 17898 32070 17910 32122
rect 17962 32070 17974 32122
rect 18026 32070 18038 32122
rect 18090 32070 18102 32122
rect 18154 32070 29110 32122
rect 29162 32070 29174 32122
rect 29226 32070 29238 32122
rect 29290 32070 29302 32122
rect 29354 32070 29366 32122
rect 29418 32070 34868 32122
rect 1104 32048 34868 32070
rect 2041 32011 2099 32017
rect 2041 31977 2053 32011
rect 2087 32008 2099 32011
rect 2958 32008 2964 32020
rect 2087 31980 2964 32008
rect 2087 31977 2099 31980
rect 2041 31971 2099 31977
rect 2958 31968 2964 31980
rect 3016 31968 3022 32020
rect 32953 32011 33011 32017
rect 32953 31977 32965 32011
rect 32999 32008 33011 32011
rect 33226 32008 33232 32020
rect 32999 31980 33232 32008
rect 32999 31977 33011 31980
rect 32953 31971 33011 31977
rect 33226 31968 33232 31980
rect 33284 31968 33290 32020
rect 33321 32011 33379 32017
rect 33321 31977 33333 32011
rect 33367 32008 33379 32011
rect 33410 32008 33416 32020
rect 33367 31980 33416 32008
rect 33367 31977 33379 31980
rect 33321 31971 33379 31977
rect 33410 31968 33416 31980
rect 33468 31968 33474 32020
rect 34241 32011 34299 32017
rect 34241 31977 34253 32011
rect 34287 32008 34299 32011
rect 35434 32008 35440 32020
rect 34287 31980 35440 32008
rect 34287 31977 34299 31980
rect 34241 31971 34299 31977
rect 35434 31968 35440 31980
rect 35492 31968 35498 32020
rect 2593 31943 2651 31949
rect 2593 31909 2605 31943
rect 2639 31940 2651 31943
rect 2774 31940 2780 31952
rect 2639 31912 2780 31940
rect 2639 31909 2651 31912
rect 2593 31903 2651 31909
rect 2774 31900 2780 31912
rect 2832 31900 2838 31952
rect 33781 31943 33839 31949
rect 33781 31909 33793 31943
rect 33827 31909 33839 31943
rect 33781 31903 33839 31909
rect 1670 31804 1676 31816
rect 1631 31776 1676 31804
rect 1670 31764 1676 31776
rect 1728 31764 1734 31816
rect 2225 31807 2283 31813
rect 2225 31773 2237 31807
rect 2271 31804 2283 31807
rect 2958 31804 2964 31816
rect 2271 31776 2964 31804
rect 2271 31773 2283 31776
rect 2225 31767 2283 31773
rect 2958 31764 2964 31776
rect 3016 31764 3022 31816
rect 32585 31807 32643 31813
rect 32585 31773 32597 31807
rect 32631 31804 32643 31807
rect 32950 31804 32956 31816
rect 32631 31776 32956 31804
rect 32631 31773 32643 31776
rect 32585 31767 32643 31773
rect 32950 31764 32956 31776
rect 33008 31764 33014 31816
rect 33594 31804 33600 31816
rect 33555 31776 33600 31804
rect 33594 31764 33600 31776
rect 33652 31764 33658 31816
rect 33796 31804 33824 31903
rect 34057 31807 34115 31813
rect 34057 31804 34069 31807
rect 33796 31776 34069 31804
rect 34057 31773 34069 31776
rect 34103 31773 34115 31807
rect 34057 31767 34115 31773
rect 1486 31668 1492 31680
rect 1447 31640 1492 31668
rect 1486 31628 1492 31640
rect 1544 31628 1550 31680
rect 1104 31578 34868 31600
rect 1104 31526 12214 31578
rect 12266 31526 12278 31578
rect 12330 31526 12342 31578
rect 12394 31526 12406 31578
rect 12458 31526 12470 31578
rect 12522 31526 23478 31578
rect 23530 31526 23542 31578
rect 23594 31526 23606 31578
rect 23658 31526 23670 31578
rect 23722 31526 23734 31578
rect 23786 31526 34868 31578
rect 1104 31504 34868 31526
rect 1394 31464 1400 31476
rect 1355 31436 1400 31464
rect 1394 31424 1400 31436
rect 1452 31424 1458 31476
rect 11882 31356 11888 31408
rect 11940 31396 11946 31408
rect 17865 31399 17923 31405
rect 17865 31396 17877 31399
rect 11940 31368 17877 31396
rect 11940 31356 11946 31368
rect 17865 31365 17877 31368
rect 17911 31365 17923 31399
rect 17865 31359 17923 31365
rect 33873 31331 33931 31337
rect 33873 31297 33885 31331
rect 33919 31328 33931 31331
rect 34330 31328 34336 31340
rect 33919 31300 34336 31328
rect 33919 31297 33931 31300
rect 33873 31291 33931 31297
rect 34330 31288 34336 31300
rect 34388 31288 34394 31340
rect 17957 31127 18015 31133
rect 17957 31093 17969 31127
rect 18003 31124 18015 31127
rect 22094 31124 22100 31136
rect 18003 31096 22100 31124
rect 18003 31093 18015 31096
rect 17957 31087 18015 31093
rect 22094 31084 22100 31096
rect 22152 31084 22158 31136
rect 33410 31124 33416 31136
rect 33371 31096 33416 31124
rect 33410 31084 33416 31096
rect 33468 31084 33474 31136
rect 33686 31084 33692 31136
rect 33744 31124 33750 31136
rect 34149 31127 34207 31133
rect 34149 31124 34161 31127
rect 33744 31096 34161 31124
rect 33744 31084 33750 31096
rect 34149 31093 34161 31096
rect 34195 31093 34207 31127
rect 34149 31087 34207 31093
rect 1104 31034 34868 31056
rect 1104 30982 6582 31034
rect 6634 30982 6646 31034
rect 6698 30982 6710 31034
rect 6762 30982 6774 31034
rect 6826 30982 6838 31034
rect 6890 30982 17846 31034
rect 17898 30982 17910 31034
rect 17962 30982 17974 31034
rect 18026 30982 18038 31034
rect 18090 30982 18102 31034
rect 18154 30982 29110 31034
rect 29162 30982 29174 31034
rect 29226 30982 29238 31034
rect 29290 30982 29302 31034
rect 29354 30982 29366 31034
rect 29418 30982 34868 31034
rect 1104 30960 34868 30982
rect 22094 30880 22100 30932
rect 22152 30920 22158 30932
rect 34054 30920 34060 30932
rect 22152 30892 34060 30920
rect 22152 30880 22158 30892
rect 34054 30880 34060 30892
rect 34112 30880 34118 30932
rect 30374 30744 30380 30796
rect 30432 30784 30438 30796
rect 34057 30787 34115 30793
rect 34057 30784 34069 30787
rect 30432 30756 34069 30784
rect 30432 30744 30438 30756
rect 34057 30753 34069 30756
rect 34103 30753 34115 30787
rect 34057 30747 34115 30753
rect 1673 30719 1731 30725
rect 1673 30685 1685 30719
rect 1719 30716 1731 30719
rect 34330 30716 34336 30728
rect 1719 30688 2084 30716
rect 34291 30688 34336 30716
rect 1719 30685 1731 30688
rect 1673 30679 1731 30685
rect 1486 30580 1492 30592
rect 1447 30552 1492 30580
rect 1486 30540 1492 30552
rect 1544 30540 1550 30592
rect 2056 30589 2084 30688
rect 34330 30676 34336 30688
rect 34388 30676 34394 30728
rect 2041 30583 2099 30589
rect 2041 30549 2053 30583
rect 2087 30580 2099 30583
rect 2130 30580 2136 30592
rect 2087 30552 2136 30580
rect 2087 30549 2099 30552
rect 2041 30543 2099 30549
rect 2130 30540 2136 30552
rect 2188 30540 2194 30592
rect 1104 30490 34868 30512
rect 1104 30438 12214 30490
rect 12266 30438 12278 30490
rect 12330 30438 12342 30490
rect 12394 30438 12406 30490
rect 12458 30438 12470 30490
rect 12522 30438 23478 30490
rect 23530 30438 23542 30490
rect 23594 30438 23606 30490
rect 23658 30438 23670 30490
rect 23722 30438 23734 30490
rect 23786 30438 34868 30490
rect 1104 30416 34868 30438
rect 33873 30379 33931 30385
rect 33873 30345 33885 30379
rect 33919 30376 33931 30379
rect 34330 30376 34336 30388
rect 33919 30348 34336 30376
rect 33919 30345 33931 30348
rect 33873 30339 33931 30345
rect 34330 30336 34336 30348
rect 34388 30336 34394 30388
rect 1949 30243 2007 30249
rect 1949 30209 1961 30243
rect 1995 30240 2007 30243
rect 33505 30243 33563 30249
rect 1995 30212 6914 30240
rect 1995 30209 2007 30212
rect 1949 30203 2007 30209
rect 2225 30175 2283 30181
rect 2225 30141 2237 30175
rect 2271 30141 2283 30175
rect 6886 30172 6914 30212
rect 33505 30209 33517 30243
rect 33551 30240 33563 30243
rect 34330 30240 34336 30252
rect 33551 30212 34336 30240
rect 33551 30209 33563 30212
rect 33505 30203 33563 30209
rect 34330 30200 34336 30212
rect 34388 30200 34394 30252
rect 18506 30172 18512 30184
rect 6886 30144 18512 30172
rect 2225 30135 2283 30141
rect 1946 30064 1952 30116
rect 2004 30104 2010 30116
rect 2240 30104 2268 30135
rect 18506 30132 18512 30144
rect 18564 30132 18570 30184
rect 2004 30076 2268 30104
rect 2004 30064 2010 30076
rect 33870 29996 33876 30048
rect 33928 30036 33934 30048
rect 34149 30039 34207 30045
rect 34149 30036 34161 30039
rect 33928 30008 34161 30036
rect 33928 29996 33934 30008
rect 34149 30005 34161 30008
rect 34195 30005 34207 30039
rect 34149 29999 34207 30005
rect 1104 29946 34868 29968
rect 1104 29894 6582 29946
rect 6634 29894 6646 29946
rect 6698 29894 6710 29946
rect 6762 29894 6774 29946
rect 6826 29894 6838 29946
rect 6890 29894 17846 29946
rect 17898 29894 17910 29946
rect 17962 29894 17974 29946
rect 18026 29894 18038 29946
rect 18090 29894 18102 29946
rect 18154 29894 29110 29946
rect 29162 29894 29174 29946
rect 29226 29894 29238 29946
rect 29290 29894 29302 29946
rect 29354 29894 29366 29946
rect 29418 29894 34868 29946
rect 1104 29872 34868 29894
rect 1946 29832 1952 29844
rect 1907 29804 1952 29832
rect 1946 29792 1952 29804
rect 2004 29792 2010 29844
rect 33594 29792 33600 29844
rect 33652 29832 33658 29844
rect 34149 29835 34207 29841
rect 34149 29832 34161 29835
rect 33652 29804 34161 29832
rect 33652 29792 33658 29804
rect 34149 29801 34161 29804
rect 34195 29801 34207 29835
rect 34149 29795 34207 29801
rect 1673 29631 1731 29637
rect 1673 29597 1685 29631
rect 1719 29628 1731 29631
rect 33873 29631 33931 29637
rect 1719 29600 2452 29628
rect 1719 29597 1731 29600
rect 1673 29591 1731 29597
rect 2424 29504 2452 29600
rect 33873 29597 33885 29631
rect 33919 29628 33931 29631
rect 34330 29628 34336 29640
rect 33919 29600 34336 29628
rect 33919 29597 33931 29600
rect 33873 29591 33931 29597
rect 34330 29588 34336 29600
rect 34388 29588 34394 29640
rect 1486 29492 1492 29504
rect 1447 29464 1492 29492
rect 1486 29452 1492 29464
rect 1544 29452 1550 29504
rect 2406 29492 2412 29504
rect 2367 29464 2412 29492
rect 2406 29452 2412 29464
rect 2464 29452 2470 29504
rect 1104 29402 34868 29424
rect 1104 29350 12214 29402
rect 12266 29350 12278 29402
rect 12330 29350 12342 29402
rect 12394 29350 12406 29402
rect 12458 29350 12470 29402
rect 12522 29350 23478 29402
rect 23530 29350 23542 29402
rect 23594 29350 23606 29402
rect 23658 29350 23670 29402
rect 23722 29350 23734 29402
rect 23786 29350 34868 29402
rect 1104 29328 34868 29350
rect 1670 29152 1676 29164
rect 1631 29124 1676 29152
rect 1670 29112 1676 29124
rect 1728 29152 1734 29164
rect 2133 29155 2191 29161
rect 2133 29152 2145 29155
rect 1728 29124 2145 29152
rect 1728 29112 1734 29124
rect 2133 29121 2145 29124
rect 2179 29121 2191 29155
rect 2133 29115 2191 29121
rect 33597 29155 33655 29161
rect 33597 29121 33609 29155
rect 33643 29152 33655 29155
rect 33870 29152 33876 29164
rect 33643 29124 33876 29152
rect 33643 29121 33655 29124
rect 33597 29115 33655 29121
rect 33870 29112 33876 29124
rect 33928 29112 33934 29164
rect 34054 29152 34060 29164
rect 34015 29124 34060 29152
rect 34054 29112 34060 29124
rect 34112 29112 34118 29164
rect 1857 29019 1915 29025
rect 1857 28985 1869 29019
rect 1903 29016 1915 29019
rect 1946 29016 1952 29028
rect 1903 28988 1952 29016
rect 1903 28985 1915 28988
rect 1857 28979 1915 28985
rect 1946 28976 1952 28988
rect 2004 28976 2010 29028
rect 34238 29016 34244 29028
rect 34199 28988 34244 29016
rect 34238 28976 34244 28988
rect 34296 28976 34302 29028
rect 33781 28951 33839 28957
rect 33781 28917 33793 28951
rect 33827 28948 33839 28951
rect 34054 28948 34060 28960
rect 33827 28920 34060 28948
rect 33827 28917 33839 28920
rect 33781 28911 33839 28917
rect 34054 28908 34060 28920
rect 34112 28908 34118 28960
rect 1104 28858 34868 28880
rect 1104 28806 6582 28858
rect 6634 28806 6646 28858
rect 6698 28806 6710 28858
rect 6762 28806 6774 28858
rect 6826 28806 6838 28858
rect 6890 28806 17846 28858
rect 17898 28806 17910 28858
rect 17962 28806 17974 28858
rect 18026 28806 18038 28858
rect 18090 28806 18102 28858
rect 18154 28806 29110 28858
rect 29162 28806 29174 28858
rect 29226 28806 29238 28858
rect 29290 28806 29302 28858
rect 29354 28806 29366 28858
rect 29418 28806 34868 28858
rect 1104 28784 34868 28806
rect 33962 28744 33968 28756
rect 33923 28716 33968 28744
rect 33962 28704 33968 28716
rect 34020 28704 34026 28756
rect 1104 28314 34868 28336
rect 1104 28262 12214 28314
rect 12266 28262 12278 28314
rect 12330 28262 12342 28314
rect 12394 28262 12406 28314
rect 12458 28262 12470 28314
rect 12522 28262 23478 28314
rect 23530 28262 23542 28314
rect 23594 28262 23606 28314
rect 23658 28262 23670 28314
rect 23722 28262 23734 28314
rect 23786 28262 34868 28314
rect 1104 28240 34868 28262
rect 20254 28200 20260 28212
rect 20215 28172 20260 28200
rect 20254 28160 20260 28172
rect 20312 28160 20318 28212
rect 1673 28067 1731 28073
rect 1673 28033 1685 28067
rect 1719 28064 1731 28067
rect 1719 28036 2084 28064
rect 1719 28033 1731 28036
rect 1673 28027 1731 28033
rect 1486 27928 1492 27940
rect 1447 27900 1492 27928
rect 1486 27888 1492 27900
rect 1544 27888 1550 27940
rect 2056 27869 2084 28036
rect 30834 28024 30840 28076
rect 30892 28064 30898 28076
rect 30929 28067 30987 28073
rect 30929 28064 30941 28067
rect 30892 28036 30941 28064
rect 30892 28024 30898 28036
rect 30929 28033 30941 28036
rect 30975 28033 30987 28067
rect 34054 28064 34060 28076
rect 34015 28036 34060 28064
rect 30929 28027 30987 28033
rect 34054 28024 34060 28036
rect 34112 28024 34118 28076
rect 34238 27928 34244 27940
rect 34199 27900 34244 27928
rect 34238 27888 34244 27900
rect 34296 27888 34302 27940
rect 2041 27863 2099 27869
rect 2041 27829 2053 27863
rect 2087 27860 2099 27863
rect 2222 27860 2228 27872
rect 2087 27832 2228 27860
rect 2087 27829 2099 27832
rect 2041 27823 2099 27829
rect 2222 27820 2228 27832
rect 2280 27820 2286 27872
rect 31113 27863 31171 27869
rect 31113 27829 31125 27863
rect 31159 27860 31171 27863
rect 34054 27860 34060 27872
rect 31159 27832 34060 27860
rect 31159 27829 31171 27832
rect 31113 27823 31171 27829
rect 34054 27820 34060 27832
rect 34112 27820 34118 27872
rect 1104 27770 34868 27792
rect 1104 27718 6582 27770
rect 6634 27718 6646 27770
rect 6698 27718 6710 27770
rect 6762 27718 6774 27770
rect 6826 27718 6838 27770
rect 6890 27718 17846 27770
rect 17898 27718 17910 27770
rect 17962 27718 17974 27770
rect 18026 27718 18038 27770
rect 18090 27718 18102 27770
rect 18154 27718 29110 27770
rect 29162 27718 29174 27770
rect 29226 27718 29238 27770
rect 29290 27718 29302 27770
rect 29354 27718 29366 27770
rect 29418 27718 34868 27770
rect 1104 27696 34868 27718
rect 19889 27591 19947 27597
rect 19889 27557 19901 27591
rect 19935 27588 19947 27591
rect 19978 27588 19984 27600
rect 19935 27560 19984 27588
rect 19935 27557 19947 27560
rect 19889 27551 19947 27557
rect 19978 27548 19984 27560
rect 20036 27548 20042 27600
rect 20901 27523 20959 27529
rect 20901 27520 20913 27523
rect 20456 27492 20913 27520
rect 6454 27412 6460 27464
rect 6512 27452 6518 27464
rect 19613 27455 19671 27461
rect 19613 27452 19625 27455
rect 6512 27424 19625 27452
rect 6512 27412 6518 27424
rect 19613 27421 19625 27424
rect 19659 27421 19671 27455
rect 19613 27415 19671 27421
rect 19797 27455 19855 27461
rect 19797 27421 19809 27455
rect 19843 27421 19855 27455
rect 19797 27415 19855 27421
rect 19981 27455 20039 27461
rect 19981 27421 19993 27455
rect 20027 27421 20039 27455
rect 19981 27415 20039 27421
rect 19812 27384 19840 27415
rect 19260 27356 19840 27384
rect 19996 27384 20024 27415
rect 20070 27412 20076 27464
rect 20128 27452 20134 27464
rect 20128 27424 20173 27452
rect 20128 27412 20134 27424
rect 20254 27412 20260 27464
rect 20312 27452 20318 27464
rect 20456 27461 20484 27492
rect 20901 27489 20913 27492
rect 20947 27489 20959 27523
rect 20901 27483 20959 27489
rect 20441 27455 20499 27461
rect 20441 27452 20453 27455
rect 20312 27424 20453 27452
rect 20312 27412 20318 27424
rect 20441 27421 20453 27424
rect 20487 27421 20499 27455
rect 20441 27415 20499 27421
rect 20622 27412 20628 27464
rect 20680 27452 20686 27464
rect 21269 27455 21327 27461
rect 21269 27452 21281 27455
rect 20680 27424 21281 27452
rect 20680 27412 20686 27424
rect 21269 27421 21281 27424
rect 21315 27421 21327 27455
rect 21269 27415 21327 27421
rect 21174 27384 21180 27396
rect 19996 27356 21180 27384
rect 18414 27276 18420 27328
rect 18472 27316 18478 27328
rect 19260 27325 19288 27356
rect 21174 27344 21180 27356
rect 21232 27344 21238 27396
rect 19245 27319 19303 27325
rect 19245 27316 19257 27319
rect 18472 27288 19257 27316
rect 18472 27276 18478 27288
rect 19245 27285 19257 27288
rect 19291 27285 19303 27319
rect 19245 27279 19303 27285
rect 20533 27319 20591 27325
rect 20533 27285 20545 27319
rect 20579 27316 20591 27319
rect 20806 27316 20812 27328
rect 20579 27288 20812 27316
rect 20579 27285 20591 27288
rect 20533 27279 20591 27285
rect 20806 27276 20812 27288
rect 20864 27276 20870 27328
rect 21634 27316 21640 27328
rect 21595 27288 21640 27316
rect 21634 27276 21640 27288
rect 21692 27276 21698 27328
rect 1104 27226 34868 27248
rect 1104 27174 12214 27226
rect 12266 27174 12278 27226
rect 12330 27174 12342 27226
rect 12394 27174 12406 27226
rect 12458 27174 12470 27226
rect 12522 27174 23478 27226
rect 23530 27174 23542 27226
rect 23594 27174 23606 27226
rect 23658 27174 23670 27226
rect 23722 27174 23734 27226
rect 23786 27174 34868 27226
rect 1104 27152 34868 27174
rect 18414 27072 18420 27124
rect 18472 27112 18478 27124
rect 18601 27115 18659 27121
rect 18601 27112 18613 27115
rect 18472 27084 18613 27112
rect 18472 27072 18478 27084
rect 18601 27081 18613 27084
rect 18647 27081 18659 27115
rect 18601 27075 18659 27081
rect 17957 26979 18015 26985
rect 17957 26945 17969 26979
rect 18003 26976 18015 26979
rect 18230 26976 18236 26988
rect 18003 26948 18236 26976
rect 18003 26945 18015 26948
rect 17957 26939 18015 26945
rect 18230 26936 18236 26948
rect 18288 26936 18294 26988
rect 18616 26976 18644 27075
rect 19334 27072 19340 27124
rect 19392 27112 19398 27124
rect 19613 27115 19671 27121
rect 19613 27112 19625 27115
rect 19392 27084 19625 27112
rect 19392 27072 19398 27084
rect 19613 27081 19625 27084
rect 19659 27081 19671 27115
rect 19613 27075 19671 27081
rect 20070 27072 20076 27124
rect 20128 27112 20134 27124
rect 21177 27115 21235 27121
rect 21177 27112 21189 27115
rect 20128 27084 21189 27112
rect 20128 27072 20134 27084
rect 21177 27081 21189 27084
rect 21223 27081 21235 27115
rect 24854 27112 24860 27124
rect 21177 27075 21235 27081
rect 22066 27084 24860 27112
rect 21634 27044 21640 27056
rect 20180 27016 21640 27044
rect 19058 26976 19064 26988
rect 18616 26948 19064 26976
rect 19058 26936 19064 26948
rect 19116 26976 19122 26988
rect 19521 26979 19579 26985
rect 19521 26976 19533 26979
rect 19116 26948 19533 26976
rect 19116 26936 19122 26948
rect 19521 26945 19533 26948
rect 19567 26945 19579 26979
rect 19886 26976 19892 26988
rect 19847 26948 19892 26976
rect 19521 26939 19579 26945
rect 16574 26800 16580 26852
rect 16632 26840 16638 26852
rect 17773 26843 17831 26849
rect 17773 26840 17785 26843
rect 16632 26812 17785 26840
rect 16632 26800 16638 26812
rect 17773 26809 17785 26812
rect 17819 26809 17831 26843
rect 19536 26840 19564 26939
rect 19886 26936 19892 26948
rect 19944 26936 19950 26988
rect 19978 26936 19984 26988
rect 20036 26976 20042 26988
rect 20073 26979 20131 26985
rect 20073 26976 20085 26979
rect 20036 26948 20085 26976
rect 20036 26936 20042 26948
rect 20073 26945 20085 26948
rect 20119 26945 20131 26979
rect 20073 26939 20131 26945
rect 20180 26840 20208 27016
rect 20254 26936 20260 26988
rect 20312 26976 20318 26988
rect 21192 26985 21220 27016
rect 21634 27004 21640 27016
rect 21692 27004 21698 27056
rect 20717 26979 20775 26985
rect 20717 26976 20729 26979
rect 20312 26948 20729 26976
rect 20312 26936 20318 26948
rect 20717 26945 20729 26948
rect 20763 26945 20775 26979
rect 20717 26939 20775 26945
rect 21177 26979 21235 26985
rect 21177 26945 21189 26979
rect 21223 26945 21235 26979
rect 21177 26939 21235 26945
rect 21361 26979 21419 26985
rect 21361 26945 21373 26979
rect 21407 26976 21419 26979
rect 21910 26976 21916 26988
rect 21407 26948 21916 26976
rect 21407 26945 21419 26948
rect 21361 26939 21419 26945
rect 21910 26936 21916 26948
rect 21968 26936 21974 26988
rect 20622 26908 20628 26920
rect 20583 26880 20628 26908
rect 20622 26868 20628 26880
rect 20680 26908 20686 26920
rect 21821 26911 21879 26917
rect 21821 26908 21833 26911
rect 20680 26880 21833 26908
rect 20680 26868 20686 26880
rect 21821 26877 21833 26880
rect 21867 26908 21879 26911
rect 22066 26908 22094 27084
rect 24854 27072 24860 27084
rect 24912 27072 24918 27124
rect 33781 26979 33839 26985
rect 33781 26945 33793 26979
rect 33827 26976 33839 26979
rect 34238 26976 34244 26988
rect 33827 26948 34244 26976
rect 33827 26945 33839 26948
rect 33781 26939 33839 26945
rect 34238 26936 34244 26948
rect 34296 26936 34302 26988
rect 21867 26880 22094 26908
rect 21867 26877 21879 26880
rect 21821 26871 21879 26877
rect 20254 26840 20260 26852
rect 19536 26812 20260 26840
rect 17773 26803 17831 26809
rect 20254 26800 20260 26812
rect 20312 26800 20318 26852
rect 18690 26732 18696 26784
rect 18748 26772 18754 26784
rect 18969 26775 19027 26781
rect 18969 26772 18981 26775
rect 18748 26744 18981 26772
rect 18748 26732 18754 26744
rect 18969 26741 18981 26744
rect 19015 26741 19027 26775
rect 20346 26772 20352 26784
rect 20307 26744 20352 26772
rect 18969 26735 19027 26741
rect 20346 26732 20352 26744
rect 20404 26732 20410 26784
rect 21910 26732 21916 26784
rect 21968 26772 21974 26784
rect 22281 26775 22339 26781
rect 22281 26772 22293 26775
rect 21968 26744 22293 26772
rect 21968 26732 21974 26744
rect 22281 26741 22293 26744
rect 22327 26772 22339 26775
rect 32306 26772 32312 26784
rect 22327 26744 32312 26772
rect 22327 26741 22339 26744
rect 22281 26735 22339 26741
rect 32306 26732 32312 26744
rect 32364 26732 32370 26784
rect 34146 26772 34152 26784
rect 34107 26744 34152 26772
rect 34146 26732 34152 26744
rect 34204 26732 34210 26784
rect 1104 26682 34868 26704
rect 1104 26630 6582 26682
rect 6634 26630 6646 26682
rect 6698 26630 6710 26682
rect 6762 26630 6774 26682
rect 6826 26630 6838 26682
rect 6890 26630 17846 26682
rect 17898 26630 17910 26682
rect 17962 26630 17974 26682
rect 18026 26630 18038 26682
rect 18090 26630 18102 26682
rect 18154 26630 29110 26682
rect 29162 26630 29174 26682
rect 29226 26630 29238 26682
rect 29290 26630 29302 26682
rect 29354 26630 29366 26682
rect 29418 26630 34868 26682
rect 1104 26608 34868 26630
rect 18230 26568 18236 26580
rect 18143 26540 18236 26568
rect 18230 26528 18236 26540
rect 18288 26568 18294 26580
rect 21082 26568 21088 26580
rect 18288 26540 21088 26568
rect 18288 26528 18294 26540
rect 21082 26528 21088 26540
rect 21140 26528 21146 26580
rect 21174 26528 21180 26580
rect 21232 26568 21238 26580
rect 21269 26571 21327 26577
rect 21269 26568 21281 26571
rect 21232 26540 21281 26568
rect 21232 26528 21238 26540
rect 21269 26537 21281 26540
rect 21315 26537 21327 26571
rect 21269 26531 21327 26537
rect 21453 26571 21511 26577
rect 21453 26537 21465 26571
rect 21499 26537 21511 26571
rect 21453 26531 21511 26537
rect 1581 26503 1639 26509
rect 1581 26469 1593 26503
rect 1627 26500 1639 26503
rect 3418 26500 3424 26512
rect 1627 26472 3424 26500
rect 1627 26469 1639 26472
rect 1581 26463 1639 26469
rect 3418 26460 3424 26472
rect 3476 26460 3482 26512
rect 18785 26503 18843 26509
rect 18785 26469 18797 26503
rect 18831 26500 18843 26503
rect 18831 26472 20024 26500
rect 18831 26469 18843 26472
rect 18785 26463 18843 26469
rect 2958 26392 2964 26444
rect 3016 26432 3022 26444
rect 19613 26435 19671 26441
rect 19613 26432 19625 26435
rect 3016 26404 19625 26432
rect 3016 26392 3022 26404
rect 19613 26401 19625 26404
rect 19659 26401 19671 26435
rect 19613 26395 19671 26401
rect 1394 26364 1400 26376
rect 1307 26336 1400 26364
rect 1394 26324 1400 26336
rect 1452 26364 1458 26376
rect 1857 26367 1915 26373
rect 1857 26364 1869 26367
rect 1452 26336 1869 26364
rect 1452 26324 1458 26336
rect 1857 26333 1869 26336
rect 1903 26333 1915 26367
rect 18690 26364 18696 26376
rect 18651 26336 18696 26364
rect 1857 26327 1915 26333
rect 18690 26324 18696 26336
rect 18748 26324 18754 26376
rect 19702 26324 19708 26376
rect 19760 26364 19766 26376
rect 19996 26373 20024 26472
rect 20346 26460 20352 26512
rect 20404 26500 20410 26512
rect 21468 26500 21496 26531
rect 20404 26472 21496 26500
rect 20404 26460 20410 26472
rect 32490 26460 32496 26512
rect 32548 26500 32554 26512
rect 34149 26503 34207 26509
rect 34149 26500 34161 26503
rect 32548 26472 34161 26500
rect 32548 26460 32554 26472
rect 34149 26469 34161 26472
rect 34195 26469 34207 26503
rect 34149 26463 34207 26469
rect 20533 26435 20591 26441
rect 20533 26432 20545 26435
rect 20088 26404 20545 26432
rect 20088 26376 20116 26404
rect 20533 26401 20545 26404
rect 20579 26401 20591 26435
rect 21910 26432 21916 26444
rect 20533 26395 20591 26401
rect 20732 26404 21916 26432
rect 19797 26367 19855 26373
rect 19797 26364 19809 26367
rect 19760 26336 19809 26364
rect 19760 26324 19766 26336
rect 19797 26333 19809 26336
rect 19843 26333 19855 26367
rect 19797 26327 19855 26333
rect 19981 26367 20039 26373
rect 19981 26333 19993 26367
rect 20027 26333 20039 26367
rect 19981 26327 20039 26333
rect 19889 26299 19947 26305
rect 19889 26265 19901 26299
rect 19935 26265 19947 26299
rect 19996 26296 20024 26327
rect 20070 26324 20076 26376
rect 20128 26364 20134 26376
rect 20128 26336 20173 26364
rect 20128 26324 20134 26336
rect 20254 26324 20260 26376
rect 20312 26364 20318 26376
rect 20732 26373 20760 26404
rect 21910 26392 21916 26404
rect 21968 26392 21974 26444
rect 20717 26367 20775 26373
rect 20312 26336 20357 26364
rect 20312 26324 20318 26336
rect 20717 26333 20729 26367
rect 20763 26333 20775 26367
rect 20717 26327 20775 26333
rect 20806 26324 20812 26376
rect 20864 26364 20870 26376
rect 20993 26367 21051 26373
rect 20993 26364 21005 26367
rect 20864 26336 21005 26364
rect 20864 26324 20870 26336
rect 20993 26333 21005 26336
rect 21039 26333 21051 26367
rect 20993 26327 21051 26333
rect 21082 26324 21088 26376
rect 21140 26364 21146 26376
rect 31294 26364 31300 26376
rect 21140 26336 31300 26364
rect 21140 26324 21146 26336
rect 31294 26324 31300 26336
rect 31352 26324 31358 26376
rect 33873 26367 33931 26373
rect 33873 26333 33885 26367
rect 33919 26364 33931 26367
rect 34330 26364 34336 26376
rect 33919 26336 34336 26364
rect 33919 26333 33931 26336
rect 33873 26327 33931 26333
rect 34330 26324 34336 26336
rect 34388 26324 34394 26376
rect 21637 26299 21695 26305
rect 21637 26296 21649 26299
rect 19996 26268 21649 26296
rect 19889 26259 19947 26265
rect 21637 26265 21649 26268
rect 21683 26265 21695 26299
rect 21637 26259 21695 26265
rect 19904 26228 19932 26259
rect 20346 26228 20352 26240
rect 19904 26200 20352 26228
rect 20346 26188 20352 26200
rect 20404 26188 20410 26240
rect 20898 26228 20904 26240
rect 20859 26200 20904 26228
rect 20898 26188 20904 26200
rect 20956 26188 20962 26240
rect 21450 26237 21456 26240
rect 21437 26231 21456 26237
rect 21437 26197 21449 26231
rect 21437 26191 21456 26197
rect 21450 26188 21456 26191
rect 21508 26188 21514 26240
rect 1104 26138 34868 26160
rect 1104 26086 12214 26138
rect 12266 26086 12278 26138
rect 12330 26086 12342 26138
rect 12394 26086 12406 26138
rect 12458 26086 12470 26138
rect 12522 26086 23478 26138
rect 23530 26086 23542 26138
rect 23594 26086 23606 26138
rect 23658 26086 23670 26138
rect 23722 26086 23734 26138
rect 23786 26086 34868 26138
rect 1104 26064 34868 26086
rect 18969 26027 19027 26033
rect 18969 25993 18981 26027
rect 19015 26024 19027 26027
rect 19058 26024 19064 26036
rect 19015 25996 19064 26024
rect 19015 25993 19027 25996
rect 18969 25987 19027 25993
rect 19058 25984 19064 25996
rect 19116 25984 19122 26036
rect 19613 26027 19671 26033
rect 19613 25993 19625 26027
rect 19659 26024 19671 26027
rect 19886 26024 19892 26036
rect 19659 25996 19892 26024
rect 19659 25993 19671 25996
rect 19613 25987 19671 25993
rect 19886 25984 19892 25996
rect 19944 25984 19950 26036
rect 20349 26027 20407 26033
rect 20349 25993 20361 26027
rect 20395 26024 20407 26027
rect 20395 25996 22094 26024
rect 20395 25993 20407 25996
rect 20349 25987 20407 25993
rect 17770 25916 17776 25968
rect 17828 25956 17834 25968
rect 17865 25959 17923 25965
rect 17865 25956 17877 25959
rect 17828 25928 17877 25956
rect 17828 25916 17834 25928
rect 17865 25925 17877 25928
rect 17911 25925 17923 25959
rect 17865 25919 17923 25925
rect 19245 25959 19303 25965
rect 19245 25925 19257 25959
rect 19291 25925 19303 25959
rect 19245 25919 19303 25925
rect 19461 25959 19519 25965
rect 19461 25925 19473 25959
rect 19507 25956 19519 25959
rect 19507 25928 20852 25956
rect 19507 25925 19519 25928
rect 19461 25919 19519 25925
rect 18601 25891 18659 25897
rect 18601 25857 18613 25891
rect 18647 25888 18659 25891
rect 18690 25888 18696 25900
rect 18647 25860 18696 25888
rect 18647 25857 18659 25860
rect 18601 25851 18659 25857
rect 18690 25848 18696 25860
rect 18748 25888 18754 25900
rect 19260 25888 19288 25919
rect 19610 25888 19616 25900
rect 18748 25860 19616 25888
rect 18748 25848 18754 25860
rect 19610 25848 19616 25860
rect 19668 25848 19674 25900
rect 19978 25848 19984 25900
rect 20036 25888 20042 25900
rect 20073 25891 20131 25897
rect 20073 25888 20085 25891
rect 20036 25860 20085 25888
rect 20036 25848 20042 25860
rect 20073 25857 20085 25860
rect 20119 25857 20131 25891
rect 20073 25851 20131 25857
rect 20254 25848 20260 25900
rect 20312 25888 20318 25900
rect 20441 25891 20499 25897
rect 20441 25888 20453 25891
rect 20312 25860 20453 25888
rect 20312 25848 20318 25860
rect 20441 25857 20453 25860
rect 20487 25857 20499 25891
rect 20441 25851 20499 25857
rect 20824 25829 20852 25928
rect 20898 25848 20904 25900
rect 20956 25888 20962 25900
rect 21269 25891 21327 25897
rect 21269 25888 21281 25891
rect 20956 25860 21281 25888
rect 20956 25848 20962 25860
rect 21269 25857 21281 25860
rect 21315 25857 21327 25891
rect 21269 25851 21327 25857
rect 19889 25823 19947 25829
rect 19889 25789 19901 25823
rect 19935 25820 19947 25823
rect 20809 25823 20867 25829
rect 19935 25792 20116 25820
rect 19935 25789 19947 25792
rect 19889 25783 19947 25789
rect 20088 25764 20116 25792
rect 20809 25789 20821 25823
rect 20855 25820 20867 25823
rect 21450 25820 21456 25832
rect 20855 25792 21456 25820
rect 20855 25789 20867 25792
rect 20809 25783 20867 25789
rect 21450 25780 21456 25792
rect 21508 25780 21514 25832
rect 22066 25820 22094 25996
rect 25130 25820 25136 25832
rect 22066 25792 25136 25820
rect 25130 25780 25136 25792
rect 25188 25780 25194 25832
rect 20070 25712 20076 25764
rect 20128 25712 20134 25764
rect 17957 25687 18015 25693
rect 17957 25653 17969 25687
rect 18003 25684 18015 25687
rect 18414 25684 18420 25696
rect 18003 25656 18420 25684
rect 18003 25653 18015 25656
rect 17957 25647 18015 25653
rect 18414 25644 18420 25656
rect 18472 25644 18478 25696
rect 19429 25687 19487 25693
rect 19429 25653 19441 25687
rect 19475 25684 19487 25687
rect 20346 25684 20352 25696
rect 19475 25656 20352 25684
rect 19475 25653 19487 25656
rect 19429 25647 19487 25653
rect 20346 25644 20352 25656
rect 20404 25644 20410 25696
rect 20990 25684 20996 25696
rect 20951 25656 20996 25684
rect 20990 25644 20996 25656
rect 21048 25684 21054 25696
rect 21821 25687 21879 25693
rect 21821 25684 21833 25687
rect 21048 25656 21833 25684
rect 21048 25644 21054 25656
rect 21821 25653 21833 25656
rect 21867 25653 21879 25687
rect 21821 25647 21879 25653
rect 1104 25594 34868 25616
rect 1104 25542 6582 25594
rect 6634 25542 6646 25594
rect 6698 25542 6710 25594
rect 6762 25542 6774 25594
rect 6826 25542 6838 25594
rect 6890 25542 17846 25594
rect 17898 25542 17910 25594
rect 17962 25542 17974 25594
rect 18026 25542 18038 25594
rect 18090 25542 18102 25594
rect 18154 25542 29110 25594
rect 29162 25542 29174 25594
rect 29226 25542 29238 25594
rect 29290 25542 29302 25594
rect 29354 25542 29366 25594
rect 29418 25542 34868 25594
rect 1104 25520 34868 25542
rect 19242 25480 19248 25492
rect 19203 25452 19248 25480
rect 19242 25440 19248 25452
rect 19300 25440 19306 25492
rect 19889 25483 19947 25489
rect 19889 25449 19901 25483
rect 19935 25480 19947 25483
rect 19978 25480 19984 25492
rect 19935 25452 19984 25480
rect 19935 25449 19947 25452
rect 19889 25443 19947 25449
rect 19978 25440 19984 25452
rect 20036 25440 20042 25492
rect 20073 25483 20131 25489
rect 20073 25449 20085 25483
rect 20119 25480 20131 25483
rect 20346 25480 20352 25492
rect 20119 25452 20352 25480
rect 20119 25449 20131 25452
rect 20073 25443 20131 25449
rect 20346 25440 20352 25452
rect 20404 25440 20410 25492
rect 18414 25372 18420 25424
rect 18472 25412 18478 25424
rect 33042 25412 33048 25424
rect 18472 25384 33048 25412
rect 18472 25372 18478 25384
rect 33042 25372 33048 25384
rect 33100 25372 33106 25424
rect 19610 25304 19616 25356
rect 19668 25344 19674 25356
rect 20346 25344 20352 25356
rect 19668 25316 20352 25344
rect 19668 25304 19674 25316
rect 20346 25304 20352 25316
rect 20404 25304 20410 25356
rect 6273 25279 6331 25285
rect 6273 25245 6285 25279
rect 6319 25276 6331 25279
rect 9122 25276 9128 25288
rect 6319 25248 9128 25276
rect 6319 25245 6331 25248
rect 6273 25239 6331 25245
rect 9122 25236 9128 25248
rect 9180 25236 9186 25288
rect 19429 25279 19487 25285
rect 19429 25245 19441 25279
rect 19475 25276 19487 25279
rect 20533 25279 20591 25285
rect 19475 25248 20484 25276
rect 19475 25245 19487 25248
rect 19429 25239 19487 25245
rect 19702 25168 19708 25220
rect 19760 25208 19766 25220
rect 20041 25211 20099 25217
rect 20041 25208 20053 25211
rect 19760 25180 20053 25208
rect 19760 25168 19766 25180
rect 20041 25177 20053 25180
rect 20087 25208 20099 25211
rect 20257 25211 20315 25217
rect 20087 25180 20208 25208
rect 20087 25177 20099 25180
rect 20041 25171 20099 25177
rect 6086 25140 6092 25152
rect 6047 25112 6092 25140
rect 6086 25100 6092 25112
rect 6144 25100 6150 25152
rect 20180 25140 20208 25180
rect 20257 25177 20269 25211
rect 20303 25208 20315 25211
rect 20346 25208 20352 25220
rect 20303 25180 20352 25208
rect 20303 25177 20315 25180
rect 20257 25171 20315 25177
rect 20346 25168 20352 25180
rect 20404 25168 20410 25220
rect 20456 25208 20484 25248
rect 20533 25245 20545 25279
rect 20579 25276 20591 25279
rect 20622 25276 20628 25288
rect 20579 25248 20628 25276
rect 20579 25245 20591 25248
rect 20533 25239 20591 25245
rect 20622 25236 20628 25248
rect 20680 25236 20686 25288
rect 20717 25279 20775 25285
rect 20717 25245 20729 25279
rect 20763 25276 20775 25279
rect 20806 25276 20812 25288
rect 20763 25248 20812 25276
rect 20763 25245 20775 25248
rect 20717 25239 20775 25245
rect 20806 25236 20812 25248
rect 20864 25236 20870 25288
rect 34054 25276 34060 25288
rect 34015 25248 34060 25276
rect 34054 25236 34060 25248
rect 34112 25236 34118 25288
rect 31846 25208 31852 25220
rect 20456 25180 31852 25208
rect 31846 25168 31852 25180
rect 31904 25168 31910 25220
rect 20625 25143 20683 25149
rect 20625 25140 20637 25143
rect 20180 25112 20637 25140
rect 20625 25109 20637 25112
rect 20671 25109 20683 25143
rect 20625 25103 20683 25109
rect 20714 25100 20720 25152
rect 20772 25140 20778 25152
rect 20990 25140 20996 25152
rect 20772 25112 20996 25140
rect 20772 25100 20778 25112
rect 20990 25100 20996 25112
rect 21048 25100 21054 25152
rect 34238 25140 34244 25152
rect 34199 25112 34244 25140
rect 34238 25100 34244 25112
rect 34296 25100 34302 25152
rect 1104 25050 34868 25072
rect 1104 24998 12214 25050
rect 12266 24998 12278 25050
rect 12330 24998 12342 25050
rect 12394 24998 12406 25050
rect 12458 24998 12470 25050
rect 12522 24998 23478 25050
rect 23530 24998 23542 25050
rect 23594 24998 23606 25050
rect 23658 24998 23670 25050
rect 23722 24998 23734 25050
rect 23786 24998 34868 25050
rect 1104 24976 34868 24998
rect 19797 24939 19855 24945
rect 19797 24905 19809 24939
rect 19843 24936 19855 24939
rect 20254 24936 20260 24948
rect 19843 24908 20260 24936
rect 19843 24905 19855 24908
rect 19797 24899 19855 24905
rect 20254 24896 20260 24908
rect 20312 24896 20318 24948
rect 1673 24803 1731 24809
rect 1673 24769 1685 24803
rect 1719 24800 1731 24803
rect 2038 24800 2044 24812
rect 1719 24772 2044 24800
rect 1719 24769 1731 24772
rect 1673 24763 1731 24769
rect 2038 24760 2044 24772
rect 2096 24760 2102 24812
rect 34054 24800 34060 24812
rect 34015 24772 34060 24800
rect 34054 24760 34060 24772
rect 34112 24760 34118 24812
rect 1486 24596 1492 24608
rect 1447 24568 1492 24596
rect 1486 24556 1492 24568
rect 1544 24556 1550 24608
rect 2038 24596 2044 24608
rect 1999 24568 2044 24596
rect 2038 24556 2044 24568
rect 2096 24556 2102 24608
rect 20438 24596 20444 24608
rect 20399 24568 20444 24596
rect 20438 24556 20444 24568
rect 20496 24556 20502 24608
rect 34238 24596 34244 24608
rect 34199 24568 34244 24596
rect 34238 24556 34244 24568
rect 34296 24556 34302 24608
rect 1104 24506 34868 24528
rect 1104 24454 6582 24506
rect 6634 24454 6646 24506
rect 6698 24454 6710 24506
rect 6762 24454 6774 24506
rect 6826 24454 6838 24506
rect 6890 24454 17846 24506
rect 17898 24454 17910 24506
rect 17962 24454 17974 24506
rect 18026 24454 18038 24506
rect 18090 24454 18102 24506
rect 18154 24454 29110 24506
rect 29162 24454 29174 24506
rect 29226 24454 29238 24506
rect 29290 24454 29302 24506
rect 29354 24454 29366 24506
rect 29418 24454 34868 24506
rect 1104 24432 34868 24454
rect 1673 24191 1731 24197
rect 1673 24157 1685 24191
rect 1719 24157 1731 24191
rect 1673 24151 1731 24157
rect 1688 24120 1716 24151
rect 2041 24123 2099 24129
rect 2041 24120 2053 24123
rect 1688 24092 2053 24120
rect 2041 24089 2053 24092
rect 2087 24120 2099 24123
rect 16574 24120 16580 24132
rect 2087 24092 16580 24120
rect 2087 24089 2099 24092
rect 2041 24083 2099 24089
rect 16574 24080 16580 24092
rect 16632 24080 16638 24132
rect 33870 24080 33876 24132
rect 33928 24120 33934 24132
rect 33965 24123 34023 24129
rect 33965 24120 33977 24123
rect 33928 24092 33977 24120
rect 33928 24080 33934 24092
rect 33965 24089 33977 24092
rect 34011 24089 34023 24123
rect 33965 24083 34023 24089
rect 34146 24080 34152 24132
rect 34204 24120 34210 24132
rect 34204 24092 34297 24120
rect 34204 24080 34210 24092
rect 1486 24052 1492 24064
rect 1447 24024 1492 24052
rect 1486 24012 1492 24024
rect 1544 24012 1550 24064
rect 20438 24012 20444 24064
rect 20496 24052 20502 24064
rect 33597 24055 33655 24061
rect 33597 24052 33609 24055
rect 20496 24024 33609 24052
rect 20496 24012 20502 24024
rect 33597 24021 33609 24024
rect 33643 24052 33655 24055
rect 34164 24052 34192 24080
rect 33643 24024 34192 24052
rect 33643 24021 33655 24024
rect 33597 24015 33655 24021
rect 1104 23962 34868 23984
rect 1104 23910 12214 23962
rect 12266 23910 12278 23962
rect 12330 23910 12342 23962
rect 12394 23910 12406 23962
rect 12458 23910 12470 23962
rect 12522 23910 23478 23962
rect 23530 23910 23542 23962
rect 23594 23910 23606 23962
rect 23658 23910 23670 23962
rect 23722 23910 23734 23962
rect 23786 23910 34868 23962
rect 1104 23888 34868 23910
rect 33781 23783 33839 23789
rect 33781 23749 33793 23783
rect 33827 23780 33839 23783
rect 34238 23780 34244 23792
rect 33827 23752 34244 23780
rect 33827 23749 33839 23752
rect 33781 23743 33839 23749
rect 34238 23740 34244 23752
rect 34296 23740 34302 23792
rect 1673 23715 1731 23721
rect 1673 23681 1685 23715
rect 1719 23712 1731 23715
rect 4062 23712 4068 23724
rect 1719 23684 4068 23712
rect 1719 23681 1731 23684
rect 1673 23675 1731 23681
rect 4062 23672 4068 23684
rect 4120 23672 4126 23724
rect 20806 23536 20812 23588
rect 20864 23576 20870 23588
rect 34057 23579 34115 23585
rect 34057 23576 34069 23579
rect 20864 23548 34069 23576
rect 20864 23536 20870 23548
rect 34057 23545 34069 23548
rect 34103 23545 34115 23579
rect 34057 23539 34115 23545
rect 1486 23508 1492 23520
rect 1447 23480 1492 23508
rect 1486 23468 1492 23480
rect 1544 23468 1550 23520
rect 1104 23418 34868 23440
rect 1104 23366 6582 23418
rect 6634 23366 6646 23418
rect 6698 23366 6710 23418
rect 6762 23366 6774 23418
rect 6826 23366 6838 23418
rect 6890 23366 17846 23418
rect 17898 23366 17910 23418
rect 17962 23366 17974 23418
rect 18026 23366 18038 23418
rect 18090 23366 18102 23418
rect 18154 23366 29110 23418
rect 29162 23366 29174 23418
rect 29226 23366 29238 23418
rect 29290 23366 29302 23418
rect 29354 23366 29366 23418
rect 29418 23366 34868 23418
rect 1104 23344 34868 23366
rect 33042 23264 33048 23316
rect 33100 23304 33106 23316
rect 33689 23307 33747 23313
rect 33689 23304 33701 23307
rect 33100 23276 33701 23304
rect 33100 23264 33106 23276
rect 33689 23273 33701 23276
rect 33735 23273 33747 23307
rect 33689 23267 33747 23273
rect 33704 23100 33732 23267
rect 34238 23236 34244 23248
rect 34199 23208 34244 23236
rect 34238 23196 34244 23208
rect 34296 23196 34302 23248
rect 34057 23103 34115 23109
rect 34057 23100 34069 23103
rect 33704 23072 34069 23100
rect 34057 23069 34069 23072
rect 34103 23069 34115 23103
rect 34057 23063 34115 23069
rect 1104 22874 34868 22896
rect 1104 22822 12214 22874
rect 12266 22822 12278 22874
rect 12330 22822 12342 22874
rect 12394 22822 12406 22874
rect 12458 22822 12470 22874
rect 12522 22822 23478 22874
rect 23530 22822 23542 22874
rect 23594 22822 23606 22874
rect 23658 22822 23670 22874
rect 23722 22822 23734 22874
rect 23786 22822 34868 22874
rect 1104 22800 34868 22822
rect 1673 22627 1731 22633
rect 1673 22593 1685 22627
rect 1719 22624 1731 22627
rect 6086 22624 6092 22636
rect 1719 22596 6092 22624
rect 1719 22593 1731 22596
rect 1673 22587 1731 22593
rect 6086 22584 6092 22596
rect 6144 22584 6150 22636
rect 18049 22627 18107 22633
rect 18049 22593 18061 22627
rect 18095 22624 18107 22627
rect 31754 22624 31760 22636
rect 18095 22596 31760 22624
rect 18095 22593 18107 22596
rect 18049 22587 18107 22593
rect 31754 22584 31760 22596
rect 31812 22584 31818 22636
rect 31846 22584 31852 22636
rect 31904 22624 31910 22636
rect 34057 22627 34115 22633
rect 34057 22624 34069 22627
rect 31904 22596 34069 22624
rect 31904 22584 31910 22596
rect 34057 22593 34069 22596
rect 34103 22593 34115 22627
rect 34057 22587 34115 22593
rect 34330 22556 34336 22568
rect 34291 22528 34336 22556
rect 34330 22516 34336 22528
rect 34388 22516 34394 22568
rect 1486 22488 1492 22500
rect 1447 22460 1492 22488
rect 1486 22448 1492 22460
rect 1544 22448 1550 22500
rect 2222 22448 2228 22500
rect 2280 22488 2286 22500
rect 17865 22491 17923 22497
rect 17865 22488 17877 22491
rect 2280 22460 17877 22488
rect 2280 22448 2286 22460
rect 17865 22457 17877 22460
rect 17911 22457 17923 22491
rect 17865 22451 17923 22457
rect 1104 22330 34868 22352
rect 1104 22278 6582 22330
rect 6634 22278 6646 22330
rect 6698 22278 6710 22330
rect 6762 22278 6774 22330
rect 6826 22278 6838 22330
rect 6890 22278 17846 22330
rect 17898 22278 17910 22330
rect 17962 22278 17974 22330
rect 18026 22278 18038 22330
rect 18090 22278 18102 22330
rect 18154 22278 29110 22330
rect 29162 22278 29174 22330
rect 29226 22278 29238 22330
rect 29290 22278 29302 22330
rect 29354 22278 29366 22330
rect 29418 22278 34868 22330
rect 1104 22256 34868 22278
rect 33965 22219 34023 22225
rect 33965 22185 33977 22219
rect 34011 22216 34023 22219
rect 34330 22216 34336 22228
rect 34011 22188 34336 22216
rect 34011 22185 34023 22188
rect 33965 22179 34023 22185
rect 34330 22176 34336 22188
rect 34388 22176 34394 22228
rect 34330 21876 34336 21888
rect 34291 21848 34336 21876
rect 34330 21836 34336 21848
rect 34388 21836 34394 21888
rect 1104 21786 34868 21808
rect 1104 21734 12214 21786
rect 12266 21734 12278 21786
rect 12330 21734 12342 21786
rect 12394 21734 12406 21786
rect 12458 21734 12470 21786
rect 12522 21734 23478 21786
rect 23530 21734 23542 21786
rect 23594 21734 23606 21786
rect 23658 21734 23670 21786
rect 23722 21734 23734 21786
rect 23786 21734 34868 21786
rect 1104 21712 34868 21734
rect 1670 21536 1676 21548
rect 1631 21508 1676 21536
rect 1670 21496 1676 21508
rect 1728 21496 1734 21548
rect 31754 21496 31760 21548
rect 31812 21536 31818 21548
rect 34057 21539 34115 21545
rect 34057 21536 34069 21539
rect 31812 21508 34069 21536
rect 31812 21496 31818 21508
rect 34057 21505 34069 21508
rect 34103 21505 34115 21539
rect 34057 21499 34115 21505
rect 34330 21468 34336 21480
rect 34291 21440 34336 21468
rect 34330 21428 34336 21440
rect 34388 21428 34394 21480
rect 1486 21332 1492 21344
rect 1447 21304 1492 21332
rect 1486 21292 1492 21304
rect 1544 21292 1550 21344
rect 1104 21242 34868 21264
rect 1104 21190 6582 21242
rect 6634 21190 6646 21242
rect 6698 21190 6710 21242
rect 6762 21190 6774 21242
rect 6826 21190 6838 21242
rect 6890 21190 17846 21242
rect 17898 21190 17910 21242
rect 17962 21190 17974 21242
rect 18026 21190 18038 21242
rect 18090 21190 18102 21242
rect 18154 21190 29110 21242
rect 29162 21190 29174 21242
rect 29226 21190 29238 21242
rect 29290 21190 29302 21242
rect 29354 21190 29366 21242
rect 29418 21190 34868 21242
rect 1104 21168 34868 21190
rect 33229 20927 33287 20933
rect 33229 20893 33241 20927
rect 33275 20924 33287 20927
rect 33502 20924 33508 20936
rect 33275 20896 33508 20924
rect 33275 20893 33287 20896
rect 33229 20887 33287 20893
rect 33502 20884 33508 20896
rect 33560 20884 33566 20936
rect 33781 20927 33839 20933
rect 33781 20893 33793 20927
rect 33827 20893 33839 20927
rect 33781 20887 33839 20893
rect 17957 20859 18015 20865
rect 17957 20825 17969 20859
rect 18003 20856 18015 20859
rect 33796 20856 33824 20887
rect 18003 20828 33824 20856
rect 18003 20825 18015 20828
rect 17957 20819 18015 20825
rect 2038 20748 2044 20800
rect 2096 20788 2102 20800
rect 17865 20791 17923 20797
rect 17865 20788 17877 20791
rect 2096 20760 17877 20788
rect 2096 20748 2102 20760
rect 17865 20757 17877 20760
rect 17911 20757 17923 20791
rect 17865 20751 17923 20757
rect 1104 20698 34868 20720
rect 1104 20646 12214 20698
rect 12266 20646 12278 20698
rect 12330 20646 12342 20698
rect 12394 20646 12406 20698
rect 12458 20646 12470 20698
rect 12522 20646 23478 20698
rect 23530 20646 23542 20698
rect 23594 20646 23606 20698
rect 23658 20646 23670 20698
rect 23722 20646 23734 20698
rect 23786 20646 34868 20698
rect 1104 20624 34868 20646
rect 33965 20587 34023 20593
rect 33965 20553 33977 20587
rect 34011 20584 34023 20587
rect 34054 20584 34060 20596
rect 34011 20556 34060 20584
rect 34011 20553 34023 20556
rect 33965 20547 34023 20553
rect 34054 20544 34060 20556
rect 34112 20544 34118 20596
rect 34146 20448 34152 20460
rect 34107 20420 34152 20448
rect 34146 20408 34152 20420
rect 34204 20408 34210 20460
rect 1394 20244 1400 20256
rect 1355 20216 1400 20244
rect 1394 20204 1400 20216
rect 1452 20204 1458 20256
rect 1104 20154 34868 20176
rect 1104 20102 6582 20154
rect 6634 20102 6646 20154
rect 6698 20102 6710 20154
rect 6762 20102 6774 20154
rect 6826 20102 6838 20154
rect 6890 20102 17846 20154
rect 17898 20102 17910 20154
rect 17962 20102 17974 20154
rect 18026 20102 18038 20154
rect 18090 20102 18102 20154
rect 18154 20102 29110 20154
rect 29162 20102 29174 20154
rect 29226 20102 29238 20154
rect 29290 20102 29302 20154
rect 29354 20102 29366 20154
rect 29418 20102 34868 20154
rect 1104 20080 34868 20102
rect 34146 20040 34152 20052
rect 34107 20012 34152 20040
rect 34146 20000 34152 20012
rect 34204 20000 34210 20052
rect 1394 19836 1400 19848
rect 1355 19808 1400 19836
rect 1394 19796 1400 19808
rect 1452 19796 1458 19848
rect 1673 19839 1731 19845
rect 1673 19805 1685 19839
rect 1719 19836 1731 19839
rect 33873 19839 33931 19845
rect 1719 19808 6914 19836
rect 1719 19805 1731 19808
rect 1673 19799 1731 19805
rect 6886 19768 6914 19808
rect 33873 19805 33885 19839
rect 33919 19836 33931 19839
rect 34330 19836 34336 19848
rect 33919 19808 34336 19836
rect 33919 19805 33931 19808
rect 33873 19799 33931 19805
rect 34330 19796 34336 19808
rect 34388 19796 34394 19848
rect 17954 19768 17960 19780
rect 6886 19740 17960 19768
rect 17954 19728 17960 19740
rect 18012 19728 18018 19780
rect 1104 19610 34868 19632
rect 1104 19558 12214 19610
rect 12266 19558 12278 19610
rect 12330 19558 12342 19610
rect 12394 19558 12406 19610
rect 12458 19558 12470 19610
rect 12522 19558 23478 19610
rect 23530 19558 23542 19610
rect 23594 19558 23606 19610
rect 23658 19558 23670 19610
rect 23722 19558 23734 19610
rect 23786 19558 34868 19610
rect 1104 19536 34868 19558
rect 1581 19499 1639 19505
rect 1581 19465 1593 19499
rect 1627 19496 1639 19499
rect 1627 19468 6914 19496
rect 1627 19465 1639 19468
rect 1581 19459 1639 19465
rect 1394 19360 1400 19372
rect 1355 19332 1400 19360
rect 1394 19320 1400 19332
rect 1452 19360 1458 19372
rect 1949 19363 2007 19369
rect 1949 19360 1961 19363
rect 1452 19332 1961 19360
rect 1452 19320 1458 19332
rect 1949 19329 1961 19332
rect 1995 19329 2007 19363
rect 6886 19360 6914 19468
rect 31754 19456 31760 19508
rect 31812 19496 31818 19508
rect 34149 19499 34207 19505
rect 34149 19496 34161 19499
rect 31812 19468 34161 19496
rect 31812 19456 31818 19468
rect 34149 19465 34161 19468
rect 34195 19465 34207 19499
rect 34149 19459 34207 19465
rect 17954 19428 17960 19440
rect 17915 19400 17960 19428
rect 17954 19388 17960 19400
rect 18012 19388 18018 19440
rect 20714 19428 20720 19440
rect 18248 19400 20720 19428
rect 18248 19360 18276 19400
rect 20714 19388 20720 19400
rect 20772 19388 20778 19440
rect 6886 19332 18276 19360
rect 1949 19323 2007 19329
rect 18322 19320 18328 19372
rect 18380 19360 18386 19372
rect 18509 19363 18567 19369
rect 18509 19360 18521 19363
rect 18380 19332 18521 19360
rect 18380 19320 18386 19332
rect 18509 19329 18521 19332
rect 18555 19360 18567 19363
rect 18969 19363 19027 19369
rect 18969 19360 18981 19363
rect 18555 19332 18981 19360
rect 18555 19329 18567 19332
rect 18509 19323 18567 19329
rect 18969 19329 18981 19332
rect 19015 19329 19027 19363
rect 18969 19323 19027 19329
rect 33873 19363 33931 19369
rect 33873 19329 33885 19363
rect 33919 19360 33931 19363
rect 34330 19360 34336 19372
rect 33919 19332 34336 19360
rect 33919 19329 33931 19332
rect 33873 19323 33931 19329
rect 34330 19320 34336 19332
rect 34388 19320 34394 19372
rect 18693 19227 18751 19233
rect 18693 19193 18705 19227
rect 18739 19224 18751 19227
rect 28718 19224 28724 19236
rect 18739 19196 28724 19224
rect 18739 19193 18751 19196
rect 18693 19187 18751 19193
rect 28718 19184 28724 19196
rect 28776 19184 28782 19236
rect 17218 19156 17224 19168
rect 17179 19128 17224 19156
rect 17218 19116 17224 19128
rect 17276 19116 17282 19168
rect 18049 19159 18107 19165
rect 18049 19125 18061 19159
rect 18095 19156 18107 19159
rect 19242 19156 19248 19168
rect 18095 19128 19248 19156
rect 18095 19125 18107 19128
rect 18049 19119 18107 19125
rect 19242 19116 19248 19128
rect 19300 19116 19306 19168
rect 1104 19066 34868 19088
rect 1104 19014 6582 19066
rect 6634 19014 6646 19066
rect 6698 19014 6710 19066
rect 6762 19014 6774 19066
rect 6826 19014 6838 19066
rect 6890 19014 17846 19066
rect 17898 19014 17910 19066
rect 17962 19014 17974 19066
rect 18026 19014 18038 19066
rect 18090 19014 18102 19066
rect 18154 19014 29110 19066
rect 29162 19014 29174 19066
rect 29226 19014 29238 19066
rect 29290 19014 29302 19066
rect 29354 19014 29366 19066
rect 29418 19014 34868 19066
rect 1104 18992 34868 19014
rect 2130 18844 2136 18896
rect 2188 18884 2194 18896
rect 29733 18887 29791 18893
rect 29733 18884 29745 18887
rect 2188 18856 29745 18884
rect 2188 18844 2194 18856
rect 29733 18853 29745 18856
rect 29779 18853 29791 18887
rect 29733 18847 29791 18853
rect 12894 18816 12900 18828
rect 1688 18788 12900 18816
rect 1688 18757 1716 18788
rect 12894 18776 12900 18788
rect 12952 18776 12958 18828
rect 17037 18819 17095 18825
rect 17037 18816 17049 18819
rect 16546 18788 17049 18816
rect 1673 18751 1731 18757
rect 1673 18717 1685 18751
rect 1719 18717 1731 18751
rect 2130 18748 2136 18760
rect 2091 18720 2136 18748
rect 1673 18711 1731 18717
rect 2130 18708 2136 18720
rect 2188 18748 2194 18760
rect 2409 18751 2467 18757
rect 2409 18748 2421 18751
rect 2188 18720 2421 18748
rect 2188 18708 2194 18720
rect 2409 18717 2421 18720
rect 2455 18717 2467 18751
rect 16546 18748 16574 18788
rect 17037 18785 17049 18788
rect 17083 18816 17095 18819
rect 17083 18788 18000 18816
rect 17083 18785 17095 18788
rect 17037 18779 17095 18785
rect 2409 18711 2467 18717
rect 6886 18720 16574 18748
rect 2314 18640 2320 18692
rect 2372 18680 2378 18692
rect 6886 18680 6914 18720
rect 17218 18708 17224 18760
rect 17276 18748 17282 18760
rect 17972 18757 18000 18788
rect 28994 18776 29000 18828
rect 29052 18816 29058 18828
rect 33410 18816 33416 18828
rect 29052 18788 33416 18816
rect 29052 18776 29058 18788
rect 33410 18776 33416 18788
rect 33468 18776 33474 18828
rect 17405 18751 17463 18757
rect 17405 18748 17417 18751
rect 17276 18720 17417 18748
rect 17276 18708 17282 18720
rect 17405 18717 17417 18720
rect 17451 18717 17463 18751
rect 17405 18711 17463 18717
rect 17957 18751 18015 18757
rect 17957 18717 17969 18751
rect 18003 18717 18015 18751
rect 17957 18711 18015 18717
rect 18601 18751 18659 18757
rect 18601 18717 18613 18751
rect 18647 18748 18659 18751
rect 18782 18748 18788 18760
rect 18647 18720 18788 18748
rect 18647 18717 18659 18720
rect 18601 18711 18659 18717
rect 18782 18708 18788 18720
rect 18840 18708 18846 18760
rect 20714 18748 20720 18760
rect 20675 18720 20720 18748
rect 20714 18708 20720 18720
rect 20772 18748 20778 18760
rect 21177 18751 21235 18757
rect 21177 18748 21189 18751
rect 20772 18720 21189 18748
rect 20772 18708 20778 18720
rect 21177 18717 21189 18720
rect 21223 18717 21235 18751
rect 21177 18711 21235 18717
rect 29178 18708 29184 18760
rect 29236 18748 29242 18760
rect 29549 18751 29607 18757
rect 29549 18748 29561 18751
rect 29236 18720 29561 18748
rect 29236 18708 29242 18720
rect 29549 18717 29561 18720
rect 29595 18717 29607 18751
rect 29549 18711 29607 18717
rect 33873 18751 33931 18757
rect 33873 18717 33885 18751
rect 33919 18748 33931 18751
rect 34330 18748 34336 18760
rect 33919 18720 34336 18748
rect 33919 18717 33931 18720
rect 33873 18711 33931 18717
rect 34330 18708 34336 18720
rect 34388 18708 34394 18760
rect 17236 18680 17264 18708
rect 2372 18652 6914 18680
rect 16546 18652 17264 18680
rect 18141 18683 18199 18689
rect 2372 18640 2378 18652
rect 1486 18612 1492 18624
rect 1447 18584 1492 18612
rect 1486 18572 1492 18584
rect 1544 18572 1550 18624
rect 1946 18612 1952 18624
rect 1907 18584 1952 18612
rect 1946 18572 1952 18584
rect 2004 18572 2010 18624
rect 2038 18572 2044 18624
rect 2096 18612 2102 18624
rect 16546 18612 16574 18652
rect 18141 18649 18153 18683
rect 18187 18680 18199 18683
rect 18230 18680 18236 18692
rect 18187 18652 18236 18680
rect 18187 18649 18199 18652
rect 18141 18643 18199 18649
rect 18230 18640 18236 18652
rect 18288 18640 18294 18692
rect 18690 18680 18696 18692
rect 18432 18652 18696 18680
rect 2096 18584 16574 18612
rect 17497 18615 17555 18621
rect 2096 18572 2102 18584
rect 17497 18581 17509 18615
rect 17543 18612 17555 18615
rect 18432 18612 18460 18652
rect 18690 18640 18696 18652
rect 18748 18640 18754 18692
rect 22094 18640 22100 18692
rect 22152 18680 22158 18692
rect 23201 18683 23259 18689
rect 23201 18680 23213 18683
rect 22152 18652 23213 18680
rect 22152 18640 22158 18652
rect 23201 18649 23213 18652
rect 23247 18649 23259 18683
rect 23201 18643 23259 18649
rect 23385 18683 23443 18689
rect 23385 18649 23397 18683
rect 23431 18680 23443 18683
rect 31754 18680 31760 18692
rect 23431 18652 31760 18680
rect 23431 18649 23443 18652
rect 23385 18643 23443 18649
rect 31754 18640 31760 18652
rect 31812 18640 31818 18692
rect 17543 18584 18460 18612
rect 18509 18615 18567 18621
rect 17543 18581 17555 18584
rect 17497 18575 17555 18581
rect 18509 18581 18521 18615
rect 18555 18612 18567 18615
rect 19058 18612 19064 18624
rect 18555 18584 19064 18612
rect 18555 18581 18567 18584
rect 18509 18575 18567 18581
rect 19058 18572 19064 18584
rect 19116 18572 19122 18624
rect 19337 18615 19395 18621
rect 19337 18581 19349 18615
rect 19383 18612 19395 18615
rect 19978 18612 19984 18624
rect 19383 18584 19984 18612
rect 19383 18581 19395 18584
rect 19337 18575 19395 18581
rect 19978 18572 19984 18584
rect 20036 18572 20042 18624
rect 20806 18612 20812 18624
rect 20767 18584 20812 18612
rect 20806 18572 20812 18584
rect 20864 18572 20870 18624
rect 29546 18572 29552 18624
rect 29604 18612 29610 18624
rect 34149 18615 34207 18621
rect 34149 18612 34161 18615
rect 29604 18584 34161 18612
rect 29604 18572 29610 18584
rect 34149 18581 34161 18584
rect 34195 18581 34207 18615
rect 34149 18575 34207 18581
rect 1104 18522 34868 18544
rect 1104 18470 12214 18522
rect 12266 18470 12278 18522
rect 12330 18470 12342 18522
rect 12394 18470 12406 18522
rect 12458 18470 12470 18522
rect 12522 18470 23478 18522
rect 23530 18470 23542 18522
rect 23594 18470 23606 18522
rect 23658 18470 23670 18522
rect 23722 18470 23734 18522
rect 23786 18470 34868 18522
rect 1104 18448 34868 18470
rect 1670 18368 1676 18420
rect 1728 18408 1734 18420
rect 2225 18411 2283 18417
rect 2225 18408 2237 18411
rect 1728 18380 2237 18408
rect 1728 18368 1734 18380
rect 2225 18377 2237 18380
rect 2271 18377 2283 18411
rect 3510 18408 3516 18420
rect 3471 18380 3516 18408
rect 2225 18371 2283 18377
rect 3510 18368 3516 18380
rect 3568 18368 3574 18420
rect 4062 18368 4068 18420
rect 4120 18408 4126 18420
rect 7101 18411 7159 18417
rect 7101 18408 7113 18411
rect 4120 18380 7113 18408
rect 4120 18368 4126 18380
rect 7101 18377 7113 18380
rect 7147 18377 7159 18411
rect 12894 18408 12900 18420
rect 12855 18380 12900 18408
rect 7101 18371 7159 18377
rect 12894 18368 12900 18380
rect 12952 18368 12958 18420
rect 16206 18408 16212 18420
rect 16167 18380 16212 18408
rect 16206 18368 16212 18380
rect 16264 18408 16270 18420
rect 17957 18411 18015 18417
rect 16264 18380 16574 18408
rect 16264 18368 16270 18380
rect 1762 18340 1768 18352
rect 1723 18312 1768 18340
rect 1762 18300 1768 18312
rect 1820 18300 1826 18352
rect 3050 18340 3056 18352
rect 3011 18312 3056 18340
rect 3050 18300 3056 18312
rect 3108 18300 3114 18352
rect 3418 18300 3424 18352
rect 3476 18340 3482 18352
rect 5537 18343 5595 18349
rect 5537 18340 5549 18343
rect 3476 18312 5549 18340
rect 3476 18300 3482 18312
rect 5537 18309 5549 18312
rect 5583 18309 5595 18343
rect 5537 18303 5595 18309
rect 6362 18300 6368 18352
rect 6420 18340 6426 18352
rect 6549 18343 6607 18349
rect 6549 18340 6561 18343
rect 6420 18312 6561 18340
rect 6420 18300 6426 18312
rect 6549 18309 6561 18312
rect 6595 18309 6607 18343
rect 6549 18303 6607 18309
rect 6914 18300 6920 18352
rect 6972 18340 6978 18352
rect 8110 18340 8116 18352
rect 6972 18312 8116 18340
rect 6972 18300 6978 18312
rect 8110 18300 8116 18312
rect 8168 18300 8174 18352
rect 16546 18340 16574 18380
rect 17957 18377 17969 18411
rect 18003 18408 18015 18411
rect 28994 18408 29000 18420
rect 18003 18380 29000 18408
rect 18003 18377 18015 18380
rect 17957 18371 18015 18377
rect 28994 18368 29000 18380
rect 29052 18368 29058 18420
rect 29178 18408 29184 18420
rect 29139 18380 29184 18408
rect 29178 18368 29184 18380
rect 29236 18368 29242 18420
rect 29914 18408 29920 18420
rect 29875 18380 29920 18408
rect 29914 18368 29920 18380
rect 29972 18368 29978 18420
rect 30006 18368 30012 18420
rect 30064 18408 30070 18420
rect 31938 18408 31944 18420
rect 30064 18380 31944 18408
rect 30064 18368 30070 18380
rect 31938 18368 31944 18380
rect 31996 18368 32002 18420
rect 17313 18343 17371 18349
rect 17313 18340 17325 18343
rect 16546 18312 17325 18340
rect 17313 18309 17325 18312
rect 17359 18309 17371 18343
rect 17313 18303 17371 18309
rect 18509 18343 18567 18349
rect 18509 18309 18521 18343
rect 18555 18340 18567 18343
rect 19978 18340 19984 18352
rect 18555 18312 19984 18340
rect 18555 18309 18567 18312
rect 18509 18303 18567 18309
rect 19978 18300 19984 18312
rect 20036 18300 20042 18352
rect 24486 18340 24492 18352
rect 24447 18312 24492 18340
rect 24486 18300 24492 18312
rect 24544 18300 24550 18352
rect 27614 18340 27620 18352
rect 27575 18312 27620 18340
rect 27614 18300 27620 18312
rect 27672 18300 27678 18352
rect 29546 18340 29552 18352
rect 29507 18312 29552 18340
rect 29546 18300 29552 18312
rect 29604 18300 29610 18352
rect 31202 18340 31208 18352
rect 31163 18312 31208 18340
rect 31202 18300 31208 18312
rect 31260 18300 31266 18352
rect 32490 18340 32496 18352
rect 32451 18312 32496 18340
rect 32490 18300 32496 18312
rect 32548 18300 32554 18352
rect 1578 18232 1584 18284
rect 1636 18272 1642 18284
rect 2409 18275 2467 18281
rect 2409 18272 2421 18275
rect 1636 18244 2421 18272
rect 1636 18232 1642 18244
rect 2409 18241 2421 18244
rect 2455 18241 2467 18275
rect 3602 18272 3608 18284
rect 3563 18244 3608 18272
rect 2409 18235 2467 18241
rect 3602 18232 3608 18244
rect 3660 18232 3666 18284
rect 6454 18232 6460 18284
rect 6512 18272 6518 18284
rect 6733 18275 6791 18281
rect 6733 18272 6745 18275
rect 6512 18244 6745 18272
rect 6512 18232 6518 18244
rect 6733 18241 6745 18244
rect 6779 18241 6791 18275
rect 7282 18272 7288 18284
rect 7243 18244 7288 18272
rect 6733 18235 6791 18241
rect 7282 18232 7288 18244
rect 7340 18232 7346 18284
rect 13081 18275 13139 18281
rect 13081 18241 13093 18275
rect 13127 18272 13139 18275
rect 15194 18272 15200 18284
rect 13127 18244 15200 18272
rect 13127 18241 13139 18244
rect 13081 18235 13139 18241
rect 15194 18232 15200 18244
rect 15252 18232 15258 18284
rect 15838 18272 15844 18284
rect 15799 18244 15844 18272
rect 15838 18232 15844 18244
rect 15896 18232 15902 18284
rect 16758 18272 16764 18284
rect 16719 18244 16764 18272
rect 16758 18232 16764 18244
rect 16816 18232 16822 18284
rect 17034 18232 17040 18284
rect 17092 18272 17098 18284
rect 17865 18275 17923 18281
rect 17865 18272 17877 18275
rect 17092 18244 17877 18272
rect 17092 18232 17098 18244
rect 17865 18241 17877 18244
rect 17911 18241 17923 18275
rect 17865 18235 17923 18241
rect 18969 18275 19027 18281
rect 18969 18241 18981 18275
rect 19015 18241 19027 18275
rect 19518 18272 19524 18284
rect 19479 18244 19524 18272
rect 18969 18235 19027 18241
rect 1854 18164 1860 18216
rect 1912 18204 1918 18216
rect 18984 18204 19012 18235
rect 19518 18232 19524 18244
rect 19576 18232 19582 18284
rect 19610 18232 19616 18284
rect 19668 18272 19674 18284
rect 19668 18244 26234 18272
rect 19668 18232 19674 18244
rect 19981 18207 20039 18213
rect 19981 18204 19993 18207
rect 1912 18176 19993 18204
rect 1912 18164 1918 18176
rect 19981 18173 19993 18176
rect 20027 18173 20039 18207
rect 19981 18167 20039 18173
rect 2406 18096 2412 18148
rect 2464 18136 2470 18148
rect 5721 18139 5779 18145
rect 2464 18108 3096 18136
rect 2464 18096 2470 18108
rect 1854 18068 1860 18080
rect 1815 18040 1860 18068
rect 1854 18028 1860 18040
rect 1912 18028 1918 18080
rect 2958 18068 2964 18080
rect 2919 18040 2964 18068
rect 2958 18028 2964 18040
rect 3016 18028 3022 18080
rect 3068 18068 3096 18108
rect 5721 18105 5733 18139
rect 5767 18136 5779 18139
rect 6914 18136 6920 18148
rect 5767 18108 6920 18136
rect 5767 18105 5779 18108
rect 5721 18099 5779 18105
rect 6914 18096 6920 18108
rect 6972 18096 6978 18148
rect 15657 18139 15715 18145
rect 15657 18136 15669 18139
rect 7024 18108 15669 18136
rect 7024 18068 7052 18108
rect 15657 18105 15669 18108
rect 15703 18105 15715 18139
rect 16942 18136 16948 18148
rect 16903 18108 16948 18136
rect 15657 18099 15715 18105
rect 16942 18096 16948 18108
rect 17000 18096 17006 18148
rect 17494 18136 17500 18148
rect 17455 18108 17500 18136
rect 17494 18096 17500 18108
rect 17552 18096 17558 18148
rect 19610 18136 19616 18148
rect 17604 18108 19616 18136
rect 3068 18040 7052 18068
rect 16758 18028 16764 18080
rect 16816 18068 16822 18080
rect 17604 18068 17632 18108
rect 19610 18096 19616 18108
rect 19668 18096 19674 18148
rect 19705 18139 19763 18145
rect 19705 18105 19717 18139
rect 19751 18136 19763 18139
rect 24673 18139 24731 18145
rect 19751 18108 22968 18136
rect 19751 18105 19763 18108
rect 19705 18099 19763 18105
rect 16816 18040 17632 18068
rect 18417 18071 18475 18077
rect 16816 18028 16822 18040
rect 18417 18037 18429 18071
rect 18463 18068 18475 18071
rect 18966 18068 18972 18080
rect 18463 18040 18972 18068
rect 18463 18037 18475 18040
rect 18417 18031 18475 18037
rect 18966 18028 18972 18040
rect 19024 18028 19030 18080
rect 19061 18071 19119 18077
rect 19061 18037 19073 18071
rect 19107 18068 19119 18071
rect 22830 18068 22836 18080
rect 19107 18040 22836 18068
rect 19107 18037 19119 18040
rect 19061 18031 19119 18037
rect 22830 18028 22836 18040
rect 22888 18028 22894 18080
rect 22940 18068 22968 18108
rect 24673 18105 24685 18139
rect 24719 18136 24731 18139
rect 25222 18136 25228 18148
rect 24719 18108 25228 18136
rect 24719 18105 24731 18108
rect 24673 18099 24731 18105
rect 25222 18096 25228 18108
rect 25280 18096 25286 18148
rect 26206 18136 26234 18244
rect 27246 18232 27252 18284
rect 27304 18272 27310 18284
rect 27433 18275 27491 18281
rect 27433 18272 27445 18275
rect 27304 18244 27445 18272
rect 27304 18232 27310 18244
rect 27433 18241 27445 18244
rect 27479 18241 27491 18275
rect 27433 18235 27491 18241
rect 29365 18275 29423 18281
rect 29365 18241 29377 18275
rect 29411 18272 29423 18275
rect 29454 18272 29460 18284
rect 29411 18244 29460 18272
rect 29411 18241 29423 18244
rect 29365 18235 29423 18241
rect 29454 18232 29460 18244
rect 29512 18232 29518 18284
rect 30009 18275 30067 18281
rect 30009 18241 30021 18275
rect 30055 18272 30067 18275
rect 30374 18272 30380 18284
rect 30055 18244 30380 18272
rect 30055 18241 30067 18244
rect 30009 18235 30067 18241
rect 30374 18232 30380 18244
rect 30432 18232 30438 18284
rect 32858 18272 32864 18284
rect 30484 18244 32864 18272
rect 30484 18136 30512 18244
rect 32858 18232 32864 18244
rect 32916 18232 32922 18284
rect 33597 18275 33655 18281
rect 33597 18241 33609 18275
rect 33643 18272 33655 18275
rect 33686 18272 33692 18284
rect 33643 18244 33692 18272
rect 33643 18241 33655 18244
rect 33597 18235 33655 18241
rect 33686 18232 33692 18244
rect 33744 18232 33750 18284
rect 34054 18272 34060 18284
rect 34015 18244 34060 18272
rect 34054 18232 34060 18244
rect 34112 18232 34118 18284
rect 26206 18108 30512 18136
rect 30926 18096 30932 18148
rect 30984 18136 30990 18148
rect 32309 18139 32367 18145
rect 32309 18136 32321 18139
rect 30984 18108 32321 18136
rect 30984 18096 30990 18108
rect 32309 18105 32321 18108
rect 32355 18105 32367 18139
rect 32309 18099 32367 18105
rect 30006 18068 30012 18080
rect 22940 18040 30012 18068
rect 30006 18028 30012 18040
rect 30064 18028 30070 18080
rect 30374 18068 30380 18080
rect 30335 18040 30380 18068
rect 30374 18028 30380 18040
rect 30432 18028 30438 18080
rect 31294 18068 31300 18080
rect 31255 18040 31300 18068
rect 31294 18028 31300 18040
rect 31352 18028 31358 18080
rect 33781 18071 33839 18077
rect 33781 18037 33793 18071
rect 33827 18068 33839 18071
rect 33962 18068 33968 18080
rect 33827 18040 33968 18068
rect 33827 18037 33839 18040
rect 33781 18031 33839 18037
rect 33962 18028 33968 18040
rect 34020 18028 34026 18080
rect 34238 18068 34244 18080
rect 34199 18040 34244 18068
rect 34238 18028 34244 18040
rect 34296 18028 34302 18080
rect 1104 17978 34868 18000
rect 1104 17926 6582 17978
rect 6634 17926 6646 17978
rect 6698 17926 6710 17978
rect 6762 17926 6774 17978
rect 6826 17926 6838 17978
rect 6890 17926 17846 17978
rect 17898 17926 17910 17978
rect 17962 17926 17974 17978
rect 18026 17926 18038 17978
rect 18090 17926 18102 17978
rect 18154 17926 29110 17978
rect 29162 17926 29174 17978
rect 29226 17926 29238 17978
rect 29290 17926 29302 17978
rect 29354 17926 29366 17978
rect 29418 17926 34868 17978
rect 1104 17904 34868 17926
rect 2590 17864 2596 17876
rect 2551 17836 2596 17864
rect 2590 17824 2596 17836
rect 2648 17824 2654 17876
rect 15838 17824 15844 17876
rect 15896 17864 15902 17876
rect 16025 17867 16083 17873
rect 16025 17864 16037 17867
rect 15896 17836 16037 17864
rect 15896 17824 15902 17836
rect 16025 17833 16037 17836
rect 16071 17864 16083 17867
rect 16669 17867 16727 17873
rect 16071 17836 16574 17864
rect 16071 17833 16083 17836
rect 16025 17827 16083 17833
rect 16546 17796 16574 17836
rect 16669 17833 16681 17867
rect 16715 17864 16727 17867
rect 16758 17864 16764 17876
rect 16715 17836 16764 17864
rect 16715 17833 16727 17836
rect 16669 17827 16727 17833
rect 16758 17824 16764 17836
rect 16816 17824 16822 17876
rect 16850 17824 16856 17876
rect 16908 17864 16914 17876
rect 17034 17864 17040 17876
rect 16908 17836 17040 17864
rect 16908 17824 16914 17836
rect 17034 17824 17040 17836
rect 17092 17824 17098 17876
rect 18509 17867 18567 17873
rect 18509 17833 18521 17867
rect 18555 17864 18567 17867
rect 18874 17864 18880 17876
rect 18555 17836 18880 17864
rect 18555 17833 18567 17836
rect 18509 17827 18567 17833
rect 18874 17824 18880 17836
rect 18932 17824 18938 17876
rect 32950 17796 32956 17808
rect 16546 17768 32956 17796
rect 32950 17756 32956 17768
rect 33008 17756 33014 17808
rect 32858 17728 32864 17740
rect 26206 17700 32864 17728
rect 1765 17663 1823 17669
rect 1765 17629 1777 17663
rect 1811 17660 1823 17663
rect 1946 17660 1952 17672
rect 1811 17632 1952 17660
rect 1811 17629 1823 17632
rect 1765 17623 1823 17629
rect 1946 17620 1952 17632
rect 2004 17620 2010 17672
rect 17402 17660 17408 17672
rect 17363 17632 17408 17660
rect 17402 17620 17408 17632
rect 17460 17620 17466 17672
rect 17957 17663 18015 17669
rect 17957 17660 17969 17663
rect 17512 17632 17969 17660
rect 2498 17592 2504 17604
rect 2459 17564 2504 17592
rect 2498 17552 2504 17564
rect 2556 17552 2562 17604
rect 8018 17552 8024 17604
rect 8076 17592 8082 17604
rect 17512 17592 17540 17632
rect 17957 17629 17969 17632
rect 18003 17629 18015 17663
rect 17957 17623 18015 17629
rect 19705 17663 19763 17669
rect 19705 17629 19717 17663
rect 19751 17660 19763 17663
rect 26206 17660 26234 17700
rect 32858 17688 32864 17700
rect 32916 17688 32922 17740
rect 19751 17632 26234 17660
rect 19751 17629 19763 17632
rect 19705 17623 19763 17629
rect 27338 17620 27344 17672
rect 27396 17660 27402 17672
rect 29825 17663 29883 17669
rect 29825 17660 29837 17663
rect 27396 17632 29837 17660
rect 27396 17620 27402 17632
rect 29825 17629 29837 17632
rect 29871 17660 29883 17663
rect 30285 17663 30343 17669
rect 30285 17660 30297 17663
rect 29871 17632 30297 17660
rect 29871 17629 29883 17632
rect 29825 17623 29883 17629
rect 30285 17629 30297 17632
rect 30331 17629 30343 17663
rect 30285 17623 30343 17629
rect 8076 17564 17540 17592
rect 17589 17595 17647 17601
rect 8076 17552 8082 17564
rect 17420 17536 17448 17564
rect 17589 17561 17601 17595
rect 17635 17592 17647 17595
rect 17770 17592 17776 17604
rect 17635 17564 17776 17592
rect 17635 17561 17647 17564
rect 17589 17555 17647 17561
rect 17770 17552 17776 17564
rect 17828 17552 17834 17604
rect 18598 17592 18604 17604
rect 18559 17564 18604 17592
rect 18598 17552 18604 17564
rect 18656 17552 18662 17604
rect 19426 17552 19432 17604
rect 19484 17592 19490 17604
rect 19521 17595 19579 17601
rect 19521 17592 19533 17595
rect 19484 17564 19533 17592
rect 19484 17552 19490 17564
rect 19521 17561 19533 17564
rect 19567 17561 19579 17595
rect 19521 17555 19579 17561
rect 30009 17595 30067 17601
rect 30009 17561 30021 17595
rect 30055 17592 30067 17595
rect 32398 17592 32404 17604
rect 30055 17564 32404 17592
rect 30055 17561 30067 17564
rect 30009 17555 30067 17561
rect 32398 17552 32404 17564
rect 32456 17552 32462 17604
rect 1857 17527 1915 17533
rect 1857 17493 1869 17527
rect 1903 17524 1915 17527
rect 2406 17524 2412 17536
rect 1903 17496 2412 17524
rect 1903 17493 1915 17496
rect 1857 17487 1915 17493
rect 2406 17484 2412 17496
rect 2464 17484 2470 17536
rect 17402 17484 17408 17536
rect 17460 17484 17466 17536
rect 18049 17527 18107 17533
rect 18049 17493 18061 17527
rect 18095 17524 18107 17527
rect 25498 17524 25504 17536
rect 18095 17496 25504 17524
rect 18095 17493 18107 17496
rect 18049 17487 18107 17493
rect 25498 17484 25504 17496
rect 25556 17484 25562 17536
rect 1104 17434 34868 17456
rect 1104 17382 12214 17434
rect 12266 17382 12278 17434
rect 12330 17382 12342 17434
rect 12394 17382 12406 17434
rect 12458 17382 12470 17434
rect 12522 17382 23478 17434
rect 23530 17382 23542 17434
rect 23594 17382 23606 17434
rect 23658 17382 23670 17434
rect 23722 17382 23734 17434
rect 23786 17382 34868 17434
rect 1104 17360 34868 17382
rect 17402 17320 17408 17332
rect 17363 17292 17408 17320
rect 17402 17280 17408 17292
rect 17460 17280 17466 17332
rect 17957 17323 18015 17329
rect 17957 17289 17969 17323
rect 18003 17320 18015 17323
rect 25866 17320 25872 17332
rect 18003 17292 25872 17320
rect 18003 17289 18015 17292
rect 17957 17283 18015 17289
rect 25866 17280 25872 17292
rect 25924 17280 25930 17332
rect 30009 17323 30067 17329
rect 30009 17289 30021 17323
rect 30055 17289 30067 17323
rect 30009 17283 30067 17289
rect 33781 17323 33839 17329
rect 33781 17289 33793 17323
rect 33827 17320 33839 17323
rect 34054 17320 34060 17332
rect 33827 17292 34060 17320
rect 33827 17289 33839 17292
rect 33781 17283 33839 17289
rect 18325 17255 18383 17261
rect 18325 17252 18337 17255
rect 6886 17224 18337 17252
rect 1673 17187 1731 17193
rect 1673 17153 1685 17187
rect 1719 17184 1731 17187
rect 6886 17184 6914 17224
rect 18325 17221 18337 17224
rect 18371 17221 18383 17255
rect 18325 17215 18383 17221
rect 18509 17255 18567 17261
rect 18509 17221 18521 17255
rect 18555 17252 18567 17255
rect 19886 17252 19892 17264
rect 18555 17224 19892 17252
rect 18555 17221 18567 17224
rect 18509 17215 18567 17221
rect 19886 17212 19892 17224
rect 19944 17212 19950 17264
rect 30024 17252 30052 17283
rect 34054 17280 34060 17292
rect 34112 17280 34118 17332
rect 30024 17224 34100 17252
rect 1719 17156 6914 17184
rect 1719 17153 1731 17156
rect 1673 17147 1731 17153
rect 17678 17144 17684 17196
rect 17736 17184 17742 17196
rect 17865 17187 17923 17193
rect 17865 17184 17877 17187
rect 17736 17156 17877 17184
rect 17736 17144 17742 17156
rect 17865 17153 17877 17156
rect 17911 17153 17923 17187
rect 17865 17147 17923 17153
rect 29454 17144 29460 17196
rect 29512 17184 29518 17196
rect 29822 17184 29828 17196
rect 29512 17156 29828 17184
rect 29512 17144 29518 17156
rect 29822 17144 29828 17156
rect 29880 17144 29886 17196
rect 33594 17184 33600 17196
rect 33555 17156 33600 17184
rect 33594 17144 33600 17156
rect 33652 17144 33658 17196
rect 34072 17193 34100 17224
rect 34057 17187 34115 17193
rect 34057 17153 34069 17187
rect 34103 17153 34115 17187
rect 34057 17147 34115 17153
rect 18598 17076 18604 17128
rect 18656 17116 18662 17128
rect 18969 17119 19027 17125
rect 18969 17116 18981 17119
rect 18656 17088 18981 17116
rect 18656 17076 18662 17088
rect 18969 17085 18981 17088
rect 19015 17116 19027 17119
rect 33134 17116 33140 17128
rect 19015 17088 33140 17116
rect 19015 17085 19027 17088
rect 18969 17079 19027 17085
rect 33134 17076 33140 17088
rect 33192 17076 33198 17128
rect 1486 17048 1492 17060
rect 1447 17020 1492 17048
rect 1486 17008 1492 17020
rect 1544 17008 1550 17060
rect 34238 17048 34244 17060
rect 34199 17020 34244 17048
rect 34238 17008 34244 17020
rect 34296 17008 34302 17060
rect 1104 16890 34868 16912
rect 1104 16838 6582 16890
rect 6634 16838 6646 16890
rect 6698 16838 6710 16890
rect 6762 16838 6774 16890
rect 6826 16838 6838 16890
rect 6890 16838 17846 16890
rect 17898 16838 17910 16890
rect 17962 16838 17974 16890
rect 18026 16838 18038 16890
rect 18090 16838 18102 16890
rect 18154 16838 29110 16890
rect 29162 16838 29174 16890
rect 29226 16838 29238 16890
rect 29290 16838 29302 16890
rect 29354 16838 29366 16890
rect 29418 16838 34868 16890
rect 1104 16816 34868 16838
rect 17678 16776 17684 16788
rect 17639 16748 17684 16776
rect 17678 16736 17684 16748
rect 17736 16736 17742 16788
rect 34330 16436 34336 16448
rect 34291 16408 34336 16436
rect 34330 16396 34336 16408
rect 34388 16396 34394 16448
rect 1104 16346 34868 16368
rect 1104 16294 12214 16346
rect 12266 16294 12278 16346
rect 12330 16294 12342 16346
rect 12394 16294 12406 16346
rect 12458 16294 12470 16346
rect 12522 16294 23478 16346
rect 23530 16294 23542 16346
rect 23594 16294 23606 16346
rect 23658 16294 23670 16346
rect 23722 16294 23734 16346
rect 23786 16294 34868 16346
rect 1104 16272 34868 16294
rect 1673 16099 1731 16105
rect 1673 16065 1685 16099
rect 1719 16096 1731 16099
rect 18506 16096 18512 16108
rect 1719 16068 18512 16096
rect 1719 16065 1731 16068
rect 1673 16059 1731 16065
rect 18506 16056 18512 16068
rect 18564 16056 18570 16108
rect 31754 15988 31760 16040
rect 31812 16028 31818 16040
rect 34057 16031 34115 16037
rect 34057 16028 34069 16031
rect 31812 16000 34069 16028
rect 31812 15988 31818 16000
rect 34057 15997 34069 16000
rect 34103 15997 34115 16031
rect 34330 16028 34336 16040
rect 34291 16000 34336 16028
rect 34057 15991 34115 15997
rect 34330 15988 34336 16000
rect 34388 15988 34394 16040
rect 1486 15892 1492 15904
rect 1447 15864 1492 15892
rect 1486 15852 1492 15864
rect 1544 15852 1550 15904
rect 1104 15802 34868 15824
rect 1104 15750 6582 15802
rect 6634 15750 6646 15802
rect 6698 15750 6710 15802
rect 6762 15750 6774 15802
rect 6826 15750 6838 15802
rect 6890 15750 17846 15802
rect 17898 15750 17910 15802
rect 17962 15750 17974 15802
rect 18026 15750 18038 15802
rect 18090 15750 18102 15802
rect 18154 15750 29110 15802
rect 29162 15750 29174 15802
rect 29226 15750 29238 15802
rect 29290 15750 29302 15802
rect 29354 15750 29366 15802
rect 29418 15750 34868 15802
rect 1104 15728 34868 15750
rect 1581 15691 1639 15697
rect 1581 15657 1593 15691
rect 1627 15688 1639 15691
rect 2498 15688 2504 15700
rect 1627 15660 2504 15688
rect 1627 15657 1639 15660
rect 1581 15651 1639 15657
rect 2498 15648 2504 15660
rect 2556 15648 2562 15700
rect 1394 15484 1400 15496
rect 1355 15456 1400 15484
rect 1394 15444 1400 15456
rect 1452 15484 1458 15496
rect 1857 15487 1915 15493
rect 1857 15484 1869 15487
rect 1452 15456 1869 15484
rect 1452 15444 1458 15456
rect 1857 15453 1869 15456
rect 1903 15453 1915 15487
rect 34054 15484 34060 15496
rect 34015 15456 34060 15484
rect 1857 15447 1915 15453
rect 34054 15444 34060 15456
rect 34112 15444 34118 15496
rect 34238 15348 34244 15360
rect 34199 15320 34244 15348
rect 34238 15308 34244 15320
rect 34296 15308 34302 15360
rect 1104 15258 34868 15280
rect 1104 15206 12214 15258
rect 12266 15206 12278 15258
rect 12330 15206 12342 15258
rect 12394 15206 12406 15258
rect 12458 15206 12470 15258
rect 12522 15206 23478 15258
rect 23530 15206 23542 15258
rect 23594 15206 23606 15258
rect 23658 15206 23670 15258
rect 23722 15206 23734 15258
rect 23786 15206 34868 15258
rect 1104 15184 34868 15206
rect 18506 15144 18512 15156
rect 18467 15116 18512 15144
rect 18506 15104 18512 15116
rect 18564 15104 18570 15156
rect 33965 15147 34023 15153
rect 33965 15113 33977 15147
rect 34011 15144 34023 15147
rect 34054 15144 34060 15156
rect 34011 15116 34060 15144
rect 34011 15113 34023 15116
rect 33965 15107 34023 15113
rect 34054 15104 34060 15116
rect 34112 15104 34118 15156
rect 18049 15079 18107 15085
rect 18049 15045 18061 15079
rect 18095 15076 18107 15079
rect 31754 15076 31760 15088
rect 18095 15048 31760 15076
rect 18095 15045 18107 15048
rect 18049 15039 18107 15045
rect 31754 15036 31760 15048
rect 31812 15036 31818 15088
rect 18601 15011 18659 15017
rect 18601 14977 18613 15011
rect 18647 15008 18659 15011
rect 18966 15008 18972 15020
rect 18647 14980 18972 15008
rect 18647 14977 18659 14980
rect 18601 14971 18659 14977
rect 18966 14968 18972 14980
rect 19024 14968 19030 15020
rect 34146 15008 34152 15020
rect 34107 14980 34152 15008
rect 34146 14968 34152 14980
rect 34204 14968 34210 15020
rect 11698 14832 11704 14884
rect 11756 14872 11762 14884
rect 17865 14875 17923 14881
rect 17865 14872 17877 14875
rect 11756 14844 17877 14872
rect 11756 14832 11762 14844
rect 17865 14841 17877 14844
rect 17911 14841 17923 14875
rect 17865 14835 17923 14841
rect 18966 14804 18972 14816
rect 18927 14776 18972 14804
rect 18966 14764 18972 14776
rect 19024 14764 19030 14816
rect 1104 14714 34868 14736
rect 1104 14662 6582 14714
rect 6634 14662 6646 14714
rect 6698 14662 6710 14714
rect 6762 14662 6774 14714
rect 6826 14662 6838 14714
rect 6890 14662 17846 14714
rect 17898 14662 17910 14714
rect 17962 14662 17974 14714
rect 18026 14662 18038 14714
rect 18090 14662 18102 14714
rect 18154 14662 29110 14714
rect 29162 14662 29174 14714
rect 29226 14662 29238 14714
rect 29290 14662 29302 14714
rect 29354 14662 29366 14714
rect 29418 14662 34868 14714
rect 1104 14640 34868 14662
rect 34146 14600 34152 14612
rect 34107 14572 34152 14600
rect 34146 14560 34152 14572
rect 34204 14560 34210 14612
rect 1673 14399 1731 14405
rect 1673 14365 1685 14399
rect 1719 14396 1731 14399
rect 11698 14396 11704 14408
rect 1719 14368 11704 14396
rect 1719 14365 1731 14368
rect 1673 14359 1731 14365
rect 11698 14356 11704 14368
rect 11756 14356 11762 14408
rect 33505 14399 33563 14405
rect 33505 14365 33517 14399
rect 33551 14396 33563 14399
rect 34330 14396 34336 14408
rect 33551 14368 34336 14396
rect 33551 14365 33563 14368
rect 33505 14359 33563 14365
rect 34330 14356 34336 14368
rect 34388 14356 34394 14408
rect 1486 14260 1492 14272
rect 1447 14232 1492 14260
rect 1486 14220 1492 14232
rect 1544 14220 1550 14272
rect 33873 14263 33931 14269
rect 33873 14229 33885 14263
rect 33919 14260 33931 14263
rect 34330 14260 34336 14272
rect 33919 14232 34336 14260
rect 33919 14229 33931 14232
rect 33873 14223 33931 14229
rect 34330 14220 34336 14232
rect 34388 14220 34394 14272
rect 1104 14170 34868 14192
rect 1104 14118 12214 14170
rect 12266 14118 12278 14170
rect 12330 14118 12342 14170
rect 12394 14118 12406 14170
rect 12458 14118 12470 14170
rect 12522 14118 23478 14170
rect 23530 14118 23542 14170
rect 23594 14118 23606 14170
rect 23658 14118 23670 14170
rect 23722 14118 23734 14170
rect 23786 14118 34868 14170
rect 1104 14096 34868 14118
rect 33134 13880 33140 13932
rect 33192 13920 33198 13932
rect 34057 13923 34115 13929
rect 34057 13920 34069 13923
rect 33192 13892 34069 13920
rect 33192 13880 33198 13892
rect 34057 13889 34069 13892
rect 34103 13889 34115 13923
rect 34057 13883 34115 13889
rect 34330 13852 34336 13864
rect 34291 13824 34336 13852
rect 34330 13812 34336 13824
rect 34388 13812 34394 13864
rect 1104 13626 34868 13648
rect 1104 13574 6582 13626
rect 6634 13574 6646 13626
rect 6698 13574 6710 13626
rect 6762 13574 6774 13626
rect 6826 13574 6838 13626
rect 6890 13574 17846 13626
rect 17898 13574 17910 13626
rect 17962 13574 17974 13626
rect 18026 13574 18038 13626
rect 18090 13574 18102 13626
rect 18154 13574 29110 13626
rect 29162 13574 29174 13626
rect 29226 13574 29238 13626
rect 29290 13574 29302 13626
rect 29354 13574 29366 13626
rect 29418 13574 34868 13626
rect 1104 13552 34868 13574
rect 34057 13311 34115 13317
rect 34057 13308 34069 13311
rect 33704 13280 34069 13308
rect 1670 13240 1676 13252
rect 1631 13212 1676 13240
rect 1670 13200 1676 13212
rect 1728 13200 1734 13252
rect 1857 13243 1915 13249
rect 1857 13209 1869 13243
rect 1903 13240 1915 13243
rect 17678 13240 17684 13252
rect 1903 13212 17684 13240
rect 1903 13209 1915 13212
rect 1857 13203 1915 13209
rect 17678 13200 17684 13212
rect 17736 13200 17742 13252
rect 1688 13172 1716 13200
rect 33704 13184 33732 13280
rect 34057 13277 34069 13280
rect 34103 13277 34115 13311
rect 34057 13271 34115 13277
rect 2133 13175 2191 13181
rect 2133 13172 2145 13175
rect 1688 13144 2145 13172
rect 2133 13141 2145 13144
rect 2179 13141 2191 13175
rect 33686 13172 33692 13184
rect 33647 13144 33692 13172
rect 2133 13135 2191 13141
rect 33686 13132 33692 13144
rect 33744 13132 33750 13184
rect 34238 13172 34244 13184
rect 34199 13144 34244 13172
rect 34238 13132 34244 13144
rect 34296 13132 34302 13184
rect 1104 13082 34868 13104
rect 1104 13030 12214 13082
rect 12266 13030 12278 13082
rect 12330 13030 12342 13082
rect 12394 13030 12406 13082
rect 12458 13030 12470 13082
rect 12522 13030 23478 13082
rect 23530 13030 23542 13082
rect 23594 13030 23606 13082
rect 23658 13030 23670 13082
rect 23722 13030 23734 13082
rect 23786 13030 34868 13082
rect 1104 13008 34868 13030
rect 1673 12835 1731 12841
rect 1673 12801 1685 12835
rect 1719 12832 1731 12835
rect 2038 12832 2044 12844
rect 1719 12804 2044 12832
rect 1719 12801 1731 12804
rect 1673 12795 1731 12801
rect 2038 12792 2044 12804
rect 2096 12792 2102 12844
rect 17770 12792 17776 12844
rect 17828 12832 17834 12844
rect 33689 12835 33747 12841
rect 33689 12832 33701 12835
rect 17828 12804 33701 12832
rect 17828 12792 17834 12804
rect 33689 12801 33701 12804
rect 33735 12832 33747 12835
rect 34057 12835 34115 12841
rect 34057 12832 34069 12835
rect 33735 12804 34069 12832
rect 33735 12801 33747 12804
rect 33689 12795 33747 12801
rect 34057 12801 34069 12804
rect 34103 12801 34115 12835
rect 34057 12795 34115 12801
rect 1486 12628 1492 12640
rect 1447 12600 1492 12628
rect 1486 12588 1492 12600
rect 1544 12588 1550 12640
rect 2038 12628 2044 12640
rect 1999 12600 2044 12628
rect 2038 12588 2044 12600
rect 2096 12588 2102 12640
rect 34238 12628 34244 12640
rect 34199 12600 34244 12628
rect 34238 12588 34244 12600
rect 34296 12588 34302 12640
rect 1104 12538 34868 12560
rect 1104 12486 6582 12538
rect 6634 12486 6646 12538
rect 6698 12486 6710 12538
rect 6762 12486 6774 12538
rect 6826 12486 6838 12538
rect 6890 12486 17846 12538
rect 17898 12486 17910 12538
rect 17962 12486 17974 12538
rect 18026 12486 18038 12538
rect 18090 12486 18102 12538
rect 18154 12486 29110 12538
rect 29162 12486 29174 12538
rect 29226 12486 29238 12538
rect 29290 12486 29302 12538
rect 29354 12486 29366 12538
rect 29418 12486 34868 12538
rect 1104 12464 34868 12486
rect 1104 11994 34868 12016
rect 1104 11942 12214 11994
rect 12266 11942 12278 11994
rect 12330 11942 12342 11994
rect 12394 11942 12406 11994
rect 12458 11942 12470 11994
rect 12522 11942 23478 11994
rect 23530 11942 23542 11994
rect 23594 11942 23606 11994
rect 23658 11942 23670 11994
rect 23722 11942 23734 11994
rect 23786 11942 34868 11994
rect 1104 11920 34868 11942
rect 17957 11747 18015 11753
rect 17957 11744 17969 11747
rect 6886 11716 17969 11744
rect 1394 11676 1400 11688
rect 1355 11648 1400 11676
rect 1394 11636 1400 11648
rect 1452 11636 1458 11688
rect 1673 11679 1731 11685
rect 1673 11645 1685 11679
rect 1719 11676 1731 11679
rect 6886 11676 6914 11716
rect 17957 11713 17969 11716
rect 18003 11713 18015 11747
rect 34057 11747 34115 11753
rect 34057 11744 34069 11747
rect 17957 11707 18015 11713
rect 26206 11716 34069 11744
rect 1719 11648 6914 11676
rect 18141 11679 18199 11685
rect 1719 11645 1731 11648
rect 1673 11639 1731 11645
rect 18141 11645 18153 11679
rect 18187 11676 18199 11679
rect 26206 11676 26234 11716
rect 34057 11713 34069 11716
rect 34103 11713 34115 11747
rect 34057 11707 34115 11713
rect 18187 11648 26234 11676
rect 18187 11645 18199 11648
rect 18141 11639 18199 11645
rect 18874 11568 18880 11620
rect 18932 11608 18938 11620
rect 19242 11608 19248 11620
rect 18932 11580 19248 11608
rect 18932 11568 18938 11580
rect 19242 11568 19248 11580
rect 19300 11568 19306 11620
rect 34238 11608 34244 11620
rect 34199 11580 34244 11608
rect 34238 11568 34244 11580
rect 34296 11568 34302 11620
rect 1104 11450 34868 11472
rect 1104 11398 6582 11450
rect 6634 11398 6646 11450
rect 6698 11398 6710 11450
rect 6762 11398 6774 11450
rect 6826 11398 6838 11450
rect 6890 11398 17846 11450
rect 17898 11398 17910 11450
rect 17962 11398 17974 11450
rect 18026 11398 18038 11450
rect 18090 11398 18102 11450
rect 18154 11398 29110 11450
rect 29162 11398 29174 11450
rect 29226 11398 29238 11450
rect 29290 11398 29302 11450
rect 29354 11398 29366 11450
rect 29418 11398 34868 11450
rect 1104 11376 34868 11398
rect 1394 11336 1400 11348
rect 1355 11308 1400 11336
rect 1394 11296 1400 11308
rect 1452 11296 1458 11348
rect 1104 10906 34868 10928
rect 1104 10854 12214 10906
rect 12266 10854 12278 10906
rect 12330 10854 12342 10906
rect 12394 10854 12406 10906
rect 12458 10854 12470 10906
rect 12522 10854 23478 10906
rect 23530 10854 23542 10906
rect 23594 10854 23606 10906
rect 23658 10854 23670 10906
rect 23722 10854 23734 10906
rect 23786 10854 34868 10906
rect 1104 10832 34868 10854
rect 1578 10792 1584 10804
rect 1539 10764 1584 10792
rect 1578 10752 1584 10764
rect 1636 10752 1642 10804
rect 1394 10656 1400 10668
rect 1355 10628 1400 10656
rect 1394 10616 1400 10628
rect 1452 10656 1458 10668
rect 1857 10659 1915 10665
rect 1857 10656 1869 10659
rect 1452 10628 1869 10656
rect 1452 10616 1458 10628
rect 1857 10625 1869 10628
rect 1903 10625 1915 10659
rect 1857 10619 1915 10625
rect 1104 10362 34868 10384
rect 1104 10310 6582 10362
rect 6634 10310 6646 10362
rect 6698 10310 6710 10362
rect 6762 10310 6774 10362
rect 6826 10310 6838 10362
rect 6890 10310 17846 10362
rect 17898 10310 17910 10362
rect 17962 10310 17974 10362
rect 18026 10310 18038 10362
rect 18090 10310 18102 10362
rect 18154 10310 29110 10362
rect 29162 10310 29174 10362
rect 29226 10310 29238 10362
rect 29290 10310 29302 10362
rect 29354 10310 29366 10362
rect 29418 10310 34868 10362
rect 1104 10288 34868 10310
rect 33594 10208 33600 10260
rect 33652 10248 33658 10260
rect 34149 10251 34207 10257
rect 34149 10248 34161 10251
rect 33652 10220 34161 10248
rect 33652 10208 33658 10220
rect 34149 10217 34161 10220
rect 34195 10217 34207 10251
rect 34149 10211 34207 10217
rect 33873 10047 33931 10053
rect 33873 10013 33885 10047
rect 33919 10044 33931 10047
rect 34330 10044 34336 10056
rect 33919 10016 34336 10044
rect 33919 10013 33931 10016
rect 33873 10007 33931 10013
rect 34330 10004 34336 10016
rect 34388 10004 34394 10056
rect 17310 9936 17316 9988
rect 17368 9976 17374 9988
rect 17405 9979 17463 9985
rect 17405 9976 17417 9979
rect 17368 9948 17417 9976
rect 17368 9936 17374 9948
rect 17405 9945 17417 9948
rect 17451 9945 17463 9979
rect 17405 9939 17463 9945
rect 17497 9911 17555 9917
rect 17497 9877 17509 9911
rect 17543 9908 17555 9911
rect 33686 9908 33692 9920
rect 17543 9880 33692 9908
rect 17543 9877 17555 9880
rect 17497 9871 17555 9877
rect 33686 9868 33692 9880
rect 33744 9868 33750 9920
rect 1104 9818 34868 9840
rect 1104 9766 12214 9818
rect 12266 9766 12278 9818
rect 12330 9766 12342 9818
rect 12394 9766 12406 9818
rect 12458 9766 12470 9818
rect 12522 9766 23478 9818
rect 23530 9766 23542 9818
rect 23594 9766 23606 9818
rect 23658 9766 23670 9818
rect 23722 9766 23734 9818
rect 23786 9766 34868 9818
rect 1104 9744 34868 9766
rect 18049 9571 18107 9577
rect 18049 9537 18061 9571
rect 18095 9568 18107 9571
rect 18506 9568 18512 9580
rect 18095 9540 18512 9568
rect 18095 9537 18107 9540
rect 18049 9531 18107 9537
rect 18506 9528 18512 9540
rect 18564 9528 18570 9580
rect 17865 9435 17923 9441
rect 17865 9432 17877 9435
rect 6886 9404 17877 9432
rect 2038 9324 2044 9376
rect 2096 9364 2102 9376
rect 6886 9364 6914 9404
rect 17865 9401 17877 9404
rect 17911 9401 17923 9435
rect 17865 9395 17923 9401
rect 18506 9364 18512 9376
rect 2096 9336 6914 9364
rect 18467 9336 18512 9364
rect 2096 9324 2102 9336
rect 18506 9324 18512 9336
rect 18564 9324 18570 9376
rect 1104 9274 34868 9296
rect 1104 9222 6582 9274
rect 6634 9222 6646 9274
rect 6698 9222 6710 9274
rect 6762 9222 6774 9274
rect 6826 9222 6838 9274
rect 6890 9222 17846 9274
rect 17898 9222 17910 9274
rect 17962 9222 17974 9274
rect 18026 9222 18038 9274
rect 18090 9222 18102 9274
rect 18154 9222 29110 9274
rect 29162 9222 29174 9274
rect 29226 9222 29238 9274
rect 29290 9222 29302 9274
rect 29354 9222 29366 9274
rect 29418 9222 34868 9274
rect 1104 9200 34868 9222
rect 1673 8959 1731 8965
rect 1673 8925 1685 8959
rect 1719 8925 1731 8959
rect 1673 8919 1731 8925
rect 1688 8888 1716 8919
rect 18230 8916 18236 8968
rect 18288 8956 18294 8968
rect 33689 8959 33747 8965
rect 33689 8956 33701 8959
rect 18288 8928 33701 8956
rect 18288 8916 18294 8928
rect 33689 8925 33701 8928
rect 33735 8956 33747 8959
rect 34057 8959 34115 8965
rect 34057 8956 34069 8959
rect 33735 8928 34069 8956
rect 33735 8925 33747 8928
rect 33689 8919 33747 8925
rect 34057 8925 34069 8928
rect 34103 8925 34115 8959
rect 34057 8919 34115 8925
rect 2041 8891 2099 8897
rect 2041 8888 2053 8891
rect 1688 8860 2053 8888
rect 2041 8857 2053 8860
rect 2087 8888 2099 8891
rect 19334 8888 19340 8900
rect 2087 8860 19340 8888
rect 2087 8857 2099 8860
rect 2041 8851 2099 8857
rect 19334 8848 19340 8860
rect 19392 8848 19398 8900
rect 1486 8820 1492 8832
rect 1447 8792 1492 8820
rect 1486 8780 1492 8792
rect 1544 8780 1550 8832
rect 34238 8820 34244 8832
rect 34199 8792 34244 8820
rect 34238 8780 34244 8792
rect 34296 8780 34302 8832
rect 1104 8730 34868 8752
rect 1104 8678 12214 8730
rect 12266 8678 12278 8730
rect 12330 8678 12342 8730
rect 12394 8678 12406 8730
rect 12458 8678 12470 8730
rect 12522 8678 23478 8730
rect 23530 8678 23542 8730
rect 23594 8678 23606 8730
rect 23658 8678 23670 8730
rect 23722 8678 23734 8730
rect 23786 8678 34868 8730
rect 1104 8656 34868 8678
rect 33781 8483 33839 8489
rect 33781 8449 33793 8483
rect 33827 8480 33839 8483
rect 34238 8480 34244 8492
rect 33827 8452 34244 8480
rect 33827 8449 33839 8452
rect 33781 8443 33839 8449
rect 34238 8440 34244 8452
rect 34296 8440 34302 8492
rect 18966 8304 18972 8356
rect 19024 8344 19030 8356
rect 34057 8347 34115 8353
rect 34057 8344 34069 8347
rect 19024 8316 34069 8344
rect 19024 8304 19030 8316
rect 34057 8313 34069 8316
rect 34103 8313 34115 8347
rect 34057 8307 34115 8313
rect 1104 8186 34868 8208
rect 1104 8134 6582 8186
rect 6634 8134 6646 8186
rect 6698 8134 6710 8186
rect 6762 8134 6774 8186
rect 6826 8134 6838 8186
rect 6890 8134 17846 8186
rect 17898 8134 17910 8186
rect 17962 8134 17974 8186
rect 18026 8134 18038 8186
rect 18090 8134 18102 8186
rect 18154 8134 29110 8186
rect 29162 8134 29174 8186
rect 29226 8134 29238 8186
rect 29290 8134 29302 8186
rect 29354 8134 29366 8186
rect 29418 8134 34868 8186
rect 1104 8112 34868 8134
rect 1673 7871 1731 7877
rect 1673 7837 1685 7871
rect 1719 7868 1731 7871
rect 10962 7868 10968 7880
rect 1719 7840 10968 7868
rect 1719 7837 1731 7840
rect 1673 7831 1731 7837
rect 10962 7828 10968 7840
rect 11020 7828 11026 7880
rect 33962 7828 33968 7880
rect 34020 7868 34026 7880
rect 34057 7871 34115 7877
rect 34057 7868 34069 7871
rect 34020 7840 34069 7868
rect 34020 7828 34026 7840
rect 34057 7837 34069 7840
rect 34103 7837 34115 7871
rect 34057 7831 34115 7837
rect 1486 7732 1492 7744
rect 1447 7704 1492 7732
rect 1486 7692 1492 7704
rect 1544 7692 1550 7744
rect 34238 7732 34244 7744
rect 34199 7704 34244 7732
rect 34238 7692 34244 7704
rect 34296 7692 34302 7744
rect 1104 7642 34868 7664
rect 1104 7590 12214 7642
rect 12266 7590 12278 7642
rect 12330 7590 12342 7642
rect 12394 7590 12406 7642
rect 12458 7590 12470 7642
rect 12522 7590 23478 7642
rect 23530 7590 23542 7642
rect 23594 7590 23606 7642
rect 23658 7590 23670 7642
rect 23722 7590 23734 7642
rect 23786 7590 34868 7642
rect 1104 7568 34868 7590
rect 1673 7395 1731 7401
rect 1673 7361 1685 7395
rect 1719 7392 1731 7395
rect 2038 7392 2044 7404
rect 1719 7364 2044 7392
rect 1719 7361 1731 7364
rect 1673 7355 1731 7361
rect 2038 7352 2044 7364
rect 2096 7352 2102 7404
rect 32398 7352 32404 7404
rect 32456 7392 32462 7404
rect 34057 7395 34115 7401
rect 34057 7392 34069 7395
rect 32456 7364 34069 7392
rect 32456 7352 32462 7364
rect 34057 7361 34069 7364
rect 34103 7361 34115 7395
rect 34057 7355 34115 7361
rect 1486 7188 1492 7200
rect 1447 7160 1492 7188
rect 1486 7148 1492 7160
rect 1544 7148 1550 7200
rect 2038 7188 2044 7200
rect 1999 7160 2044 7188
rect 2038 7148 2044 7160
rect 2096 7148 2102 7200
rect 34238 7188 34244 7200
rect 34199 7160 34244 7188
rect 34238 7148 34244 7160
rect 34296 7148 34302 7200
rect 1104 7098 34868 7120
rect 1104 7046 6582 7098
rect 6634 7046 6646 7098
rect 6698 7046 6710 7098
rect 6762 7046 6774 7098
rect 6826 7046 6838 7098
rect 6890 7046 17846 7098
rect 17898 7046 17910 7098
rect 17962 7046 17974 7098
rect 18026 7046 18038 7098
rect 18090 7046 18102 7098
rect 18154 7046 29110 7098
rect 29162 7046 29174 7098
rect 29226 7046 29238 7098
rect 29290 7046 29302 7098
rect 29354 7046 29366 7098
rect 29418 7046 34868 7098
rect 1104 7024 34868 7046
rect 1104 6554 34868 6576
rect 1104 6502 12214 6554
rect 12266 6502 12278 6554
rect 12330 6502 12342 6554
rect 12394 6502 12406 6554
rect 12458 6502 12470 6554
rect 12522 6502 23478 6554
rect 23530 6502 23542 6554
rect 23594 6502 23606 6554
rect 23658 6502 23670 6554
rect 23722 6502 23734 6554
rect 23786 6502 34868 6554
rect 1104 6480 34868 6502
rect 1673 6307 1731 6313
rect 1673 6273 1685 6307
rect 1719 6304 1731 6307
rect 2958 6304 2964 6316
rect 1719 6276 2964 6304
rect 1719 6273 1731 6276
rect 1673 6267 1731 6273
rect 2958 6264 2964 6276
rect 3016 6264 3022 6316
rect 33781 6307 33839 6313
rect 33781 6273 33793 6307
rect 33827 6304 33839 6307
rect 34238 6304 34244 6316
rect 33827 6276 34244 6304
rect 33827 6273 33839 6276
rect 33781 6267 33839 6273
rect 34238 6264 34244 6276
rect 34296 6264 34302 6316
rect 1486 6168 1492 6180
rect 1447 6140 1492 6168
rect 1486 6128 1492 6140
rect 1544 6128 1550 6180
rect 34057 6171 34115 6177
rect 34057 6168 34069 6171
rect 26206 6140 34069 6168
rect 19978 6060 19984 6112
rect 20036 6100 20042 6112
rect 26206 6100 26234 6140
rect 34057 6137 34069 6140
rect 34103 6137 34115 6171
rect 34057 6131 34115 6137
rect 20036 6072 26234 6100
rect 20036 6060 20042 6072
rect 1104 6010 34868 6032
rect 1104 5958 6582 6010
rect 6634 5958 6646 6010
rect 6698 5958 6710 6010
rect 6762 5958 6774 6010
rect 6826 5958 6838 6010
rect 6890 5958 17846 6010
rect 17898 5958 17910 6010
rect 17962 5958 17974 6010
rect 18026 5958 18038 6010
rect 18090 5958 18102 6010
rect 18154 5958 29110 6010
rect 29162 5958 29174 6010
rect 29226 5958 29238 6010
rect 29290 5958 29302 6010
rect 29354 5958 29366 6010
rect 29418 5958 34868 6010
rect 1104 5936 34868 5958
rect 34330 5556 34336 5568
rect 34291 5528 34336 5556
rect 34330 5516 34336 5528
rect 34388 5516 34394 5568
rect 1104 5466 34868 5488
rect 1104 5414 12214 5466
rect 12266 5414 12278 5466
rect 12330 5414 12342 5466
rect 12394 5414 12406 5466
rect 12458 5414 12470 5466
rect 12522 5414 23478 5466
rect 23530 5414 23542 5466
rect 23594 5414 23606 5466
rect 23658 5414 23670 5466
rect 23722 5414 23734 5466
rect 23786 5414 34868 5466
rect 1104 5392 34868 5414
rect 10962 5352 10968 5364
rect 10923 5324 10968 5352
rect 10962 5312 10968 5324
rect 11020 5312 11026 5364
rect 1673 5219 1731 5225
rect 1673 5185 1685 5219
rect 1719 5216 1731 5219
rect 11149 5219 11207 5225
rect 1719 5188 6914 5216
rect 1719 5185 1731 5188
rect 1673 5179 1731 5185
rect 6886 5148 6914 5188
rect 11149 5185 11161 5219
rect 11195 5216 11207 5219
rect 13630 5216 13636 5228
rect 11195 5188 13636 5216
rect 11195 5185 11207 5188
rect 11149 5179 11207 5185
rect 13630 5176 13636 5188
rect 13688 5176 13694 5228
rect 17770 5148 17776 5160
rect 6886 5120 17776 5148
rect 17770 5108 17776 5120
rect 17828 5108 17834 5160
rect 30098 5108 30104 5160
rect 30156 5148 30162 5160
rect 34057 5151 34115 5157
rect 34057 5148 34069 5151
rect 30156 5120 34069 5148
rect 30156 5108 30162 5120
rect 34057 5117 34069 5120
rect 34103 5117 34115 5151
rect 34330 5148 34336 5160
rect 34291 5120 34336 5148
rect 34057 5111 34115 5117
rect 34330 5108 34336 5120
rect 34388 5108 34394 5160
rect 1486 5012 1492 5024
rect 1447 4984 1492 5012
rect 1486 4972 1492 4984
rect 1544 4972 1550 5024
rect 1104 4922 34868 4944
rect 1104 4870 6582 4922
rect 6634 4870 6646 4922
rect 6698 4870 6710 4922
rect 6762 4870 6774 4922
rect 6826 4870 6838 4922
rect 6890 4870 17846 4922
rect 17898 4870 17910 4922
rect 17962 4870 17974 4922
rect 18026 4870 18038 4922
rect 18090 4870 18102 4922
rect 18154 4870 29110 4922
rect 29162 4870 29174 4922
rect 29226 4870 29238 4922
rect 29290 4870 29302 4922
rect 29354 4870 29366 4922
rect 29418 4870 34868 4922
rect 1104 4848 34868 4870
rect 17770 4700 17776 4752
rect 17828 4740 17834 4752
rect 17865 4743 17923 4749
rect 17865 4740 17877 4743
rect 17828 4712 17877 4740
rect 17828 4700 17834 4712
rect 17865 4709 17877 4712
rect 17911 4709 17923 4743
rect 17865 4703 17923 4709
rect 30098 4672 30104 4684
rect 18524 4644 30104 4672
rect 18417 4607 18475 4613
rect 18417 4604 18429 4607
rect 6886 4576 18429 4604
rect 1394 4468 1400 4480
rect 1355 4440 1400 4468
rect 1394 4428 1400 4440
rect 1452 4428 1458 4480
rect 2038 4428 2044 4480
rect 2096 4468 2102 4480
rect 6886 4468 6914 4576
rect 18417 4573 18429 4576
rect 18463 4573 18475 4607
rect 18417 4567 18475 4573
rect 18049 4539 18107 4545
rect 18049 4505 18061 4539
rect 18095 4536 18107 4539
rect 18524 4536 18552 4644
rect 30098 4632 30104 4644
rect 30156 4632 30162 4684
rect 34057 4607 34115 4613
rect 34057 4604 34069 4607
rect 33704 4576 34069 4604
rect 18095 4508 18552 4536
rect 18601 4539 18659 4545
rect 18095 4505 18107 4508
rect 18049 4499 18107 4505
rect 18601 4505 18613 4539
rect 18647 4536 18659 4539
rect 20346 4536 20352 4548
rect 18647 4508 20352 4536
rect 18647 4505 18659 4508
rect 18601 4499 18659 4505
rect 20346 4496 20352 4508
rect 20404 4496 20410 4548
rect 2096 4440 6914 4468
rect 2096 4428 2102 4440
rect 17586 4428 17592 4480
rect 17644 4468 17650 4480
rect 33704 4477 33732 4576
rect 34057 4573 34069 4576
rect 34103 4573 34115 4607
rect 34057 4567 34115 4573
rect 33689 4471 33747 4477
rect 33689 4468 33701 4471
rect 17644 4440 33701 4468
rect 17644 4428 17650 4440
rect 33689 4437 33701 4440
rect 33735 4437 33747 4471
rect 34238 4468 34244 4480
rect 34199 4440 34244 4468
rect 33689 4431 33747 4437
rect 34238 4428 34244 4440
rect 34296 4428 34302 4480
rect 1104 4378 34868 4400
rect 1104 4326 12214 4378
rect 12266 4326 12278 4378
rect 12330 4326 12342 4378
rect 12394 4326 12406 4378
rect 12458 4326 12470 4378
rect 12522 4326 23478 4378
rect 23530 4326 23542 4378
rect 23594 4326 23606 4378
rect 23658 4326 23670 4378
rect 23722 4326 23734 4378
rect 23786 4326 34868 4378
rect 1104 4304 34868 4326
rect 1394 4128 1400 4140
rect 1355 4100 1400 4128
rect 1394 4088 1400 4100
rect 1452 4088 1458 4140
rect 1857 4131 1915 4137
rect 1857 4097 1869 4131
rect 1903 4128 1915 4131
rect 3050 4128 3056 4140
rect 1903 4100 3056 4128
rect 1903 4097 1915 4100
rect 1857 4091 1915 4097
rect 3050 4088 3056 4100
rect 3108 4088 3114 4140
rect 33413 4131 33471 4137
rect 33413 4097 33425 4131
rect 33459 4128 33471 4131
rect 33870 4128 33876 4140
rect 33459 4100 33876 4128
rect 33459 4097 33471 4100
rect 33413 4091 33471 4097
rect 33870 4088 33876 4100
rect 33928 4128 33934 4140
rect 34057 4131 34115 4137
rect 34057 4128 34069 4131
rect 33928 4100 34069 4128
rect 33928 4088 33934 4100
rect 34057 4097 34069 4100
rect 34103 4097 34115 4131
rect 34057 4091 34115 4097
rect 1581 3995 1639 4001
rect 1581 3961 1593 3995
rect 1627 3992 1639 3995
rect 11606 3992 11612 4004
rect 1627 3964 11612 3992
rect 1627 3961 1639 3964
rect 1581 3955 1639 3961
rect 11606 3952 11612 3964
rect 11664 3952 11670 4004
rect 2038 3924 2044 3936
rect 1999 3896 2044 3924
rect 2038 3884 2044 3896
rect 2096 3884 2102 3936
rect 2317 3927 2375 3933
rect 2317 3893 2329 3927
rect 2363 3924 2375 3927
rect 3050 3924 3056 3936
rect 2363 3896 3056 3924
rect 2363 3893 2375 3896
rect 2317 3887 2375 3893
rect 3050 3884 3056 3896
rect 3108 3884 3114 3936
rect 33781 3927 33839 3933
rect 33781 3893 33793 3927
rect 33827 3924 33839 3927
rect 33870 3924 33876 3936
rect 33827 3896 33876 3924
rect 33827 3893 33839 3896
rect 33781 3887 33839 3893
rect 33870 3884 33876 3896
rect 33928 3884 33934 3936
rect 34238 3924 34244 3936
rect 34199 3896 34244 3924
rect 34238 3884 34244 3896
rect 34296 3884 34302 3936
rect 1104 3834 34868 3856
rect 1104 3782 6582 3834
rect 6634 3782 6646 3834
rect 6698 3782 6710 3834
rect 6762 3782 6774 3834
rect 6826 3782 6838 3834
rect 6890 3782 17846 3834
rect 17898 3782 17910 3834
rect 17962 3782 17974 3834
rect 18026 3782 18038 3834
rect 18090 3782 18102 3834
rect 18154 3782 29110 3834
rect 29162 3782 29174 3834
rect 29226 3782 29238 3834
rect 29290 3782 29302 3834
rect 29354 3782 29366 3834
rect 29418 3782 34868 3834
rect 1104 3760 34868 3782
rect 8110 3720 8116 3732
rect 8071 3692 8116 3720
rect 8110 3680 8116 3692
rect 8168 3680 8174 3732
rect 14550 3680 14556 3732
rect 14608 3720 14614 3732
rect 18325 3723 18383 3729
rect 18325 3720 18337 3723
rect 14608 3692 18337 3720
rect 14608 3680 14614 3692
rect 18325 3689 18337 3692
rect 18371 3689 18383 3723
rect 20530 3720 20536 3732
rect 18325 3683 18383 3689
rect 18432 3692 20536 3720
rect 14 3612 20 3664
rect 72 3652 78 3664
rect 2133 3655 2191 3661
rect 2133 3652 2145 3655
rect 72 3624 2145 3652
rect 72 3612 78 3624
rect 2133 3621 2145 3624
rect 2179 3621 2191 3655
rect 2133 3615 2191 3621
rect 2501 3655 2559 3661
rect 2501 3621 2513 3655
rect 2547 3621 2559 3655
rect 2501 3615 2559 3621
rect 2516 3584 2544 3615
rect 6822 3612 6828 3664
rect 6880 3652 6886 3664
rect 13722 3652 13728 3664
rect 6880 3624 13728 3652
rect 6880 3612 6886 3624
rect 13722 3612 13728 3624
rect 13780 3612 13786 3664
rect 17402 3652 17408 3664
rect 16546 3624 17408 3652
rect 1688 3556 2544 3584
rect 1688 3525 1716 3556
rect 4430 3544 4436 3596
rect 4488 3584 4494 3596
rect 16546 3584 16574 3624
rect 17402 3612 17408 3624
rect 17460 3612 17466 3664
rect 18049 3655 18107 3661
rect 18049 3621 18061 3655
rect 18095 3652 18107 3655
rect 18432 3652 18460 3692
rect 20530 3680 20536 3692
rect 20588 3680 20594 3732
rect 32861 3723 32919 3729
rect 32861 3689 32873 3723
rect 32907 3720 32919 3723
rect 34514 3720 34520 3732
rect 32907 3692 34520 3720
rect 32907 3689 32919 3692
rect 32861 3683 32919 3689
rect 34514 3680 34520 3692
rect 34572 3680 34578 3732
rect 18095 3624 18460 3652
rect 18095 3621 18107 3624
rect 18049 3615 18107 3621
rect 18506 3612 18512 3664
rect 18564 3652 18570 3664
rect 33689 3655 33747 3661
rect 18564 3624 30236 3652
rect 18564 3612 18570 3624
rect 4488 3556 16574 3584
rect 4488 3544 4494 3556
rect 17126 3544 17132 3596
rect 17184 3584 17190 3596
rect 30208 3584 30236 3624
rect 33689 3621 33701 3655
rect 33735 3652 33747 3655
rect 34790 3652 34796 3664
rect 33735 3624 34796 3652
rect 33735 3621 33747 3624
rect 33689 3615 33747 3621
rect 34790 3612 34796 3624
rect 34848 3612 34854 3664
rect 34057 3587 34115 3593
rect 34057 3584 34069 3587
rect 17184 3556 30052 3584
rect 30208 3556 34069 3584
rect 17184 3544 17190 3556
rect 1673 3519 1731 3525
rect 1673 3485 1685 3519
rect 1719 3485 1731 3519
rect 1673 3479 1731 3485
rect 1854 3476 1860 3528
rect 1912 3516 1918 3528
rect 1949 3519 2007 3525
rect 1949 3516 1961 3519
rect 1912 3488 1961 3516
rect 1912 3476 1918 3488
rect 1949 3485 1961 3488
rect 1995 3485 2007 3519
rect 1949 3479 2007 3485
rect 2038 3476 2044 3528
rect 2096 3516 2102 3528
rect 2685 3519 2743 3525
rect 2685 3516 2697 3519
rect 2096 3488 2697 3516
rect 2096 3476 2102 3488
rect 2685 3485 2697 3488
rect 2731 3485 2743 3519
rect 16666 3516 16672 3528
rect 16627 3488 16672 3516
rect 2685 3479 2743 3485
rect 16666 3476 16672 3488
rect 16724 3476 16730 3528
rect 17218 3476 17224 3528
rect 17276 3516 17282 3528
rect 17865 3519 17923 3525
rect 17865 3516 17877 3519
rect 17276 3488 17877 3516
rect 17276 3476 17282 3488
rect 17865 3485 17877 3488
rect 17911 3485 17923 3519
rect 17865 3479 17923 3485
rect 18509 3519 18567 3525
rect 18509 3485 18521 3519
rect 18555 3516 18567 3519
rect 29730 3516 29736 3528
rect 18555 3488 29736 3516
rect 18555 3485 18567 3488
rect 18509 3479 18567 3485
rect 29730 3476 29736 3488
rect 29788 3476 29794 3528
rect 30024 3516 30052 3556
rect 34057 3553 34069 3556
rect 34103 3553 34115 3587
rect 34057 3547 34115 3553
rect 31846 3516 31852 3528
rect 30024 3488 31852 3516
rect 31846 3476 31852 3488
rect 31904 3476 31910 3528
rect 32398 3516 32404 3528
rect 32359 3488 32404 3516
rect 32398 3476 32404 3488
rect 32456 3476 32462 3528
rect 33493 3519 33551 3525
rect 33493 3516 33505 3519
rect 32508 3488 33505 3516
rect 4246 3408 4252 3460
rect 4304 3448 4310 3460
rect 17770 3448 17776 3460
rect 4304 3420 17776 3448
rect 4304 3408 4310 3420
rect 17770 3408 17776 3420
rect 17828 3408 17834 3460
rect 19150 3408 19156 3460
rect 19208 3448 19214 3460
rect 19613 3451 19671 3457
rect 19613 3448 19625 3451
rect 19208 3420 19625 3448
rect 19208 3408 19214 3420
rect 19613 3417 19625 3420
rect 19659 3417 19671 3451
rect 19613 3411 19671 3417
rect 19702 3408 19708 3460
rect 19760 3448 19766 3460
rect 32508 3448 32536 3488
rect 33493 3485 33505 3488
rect 33539 3485 33551 3519
rect 33493 3479 33551 3485
rect 19760 3420 32536 3448
rect 34241 3451 34299 3457
rect 19760 3408 19766 3420
rect 34241 3417 34253 3451
rect 34287 3448 34299 3451
rect 34514 3448 34520 3460
rect 34287 3420 34520 3448
rect 34287 3417 34299 3420
rect 34241 3411 34299 3417
rect 34514 3408 34520 3420
rect 34572 3448 34578 3460
rect 35434 3448 35440 3460
rect 34572 3420 35440 3448
rect 34572 3408 34578 3420
rect 35434 3408 35440 3420
rect 35492 3408 35498 3460
rect 658 3340 664 3392
rect 716 3380 722 3392
rect 1489 3383 1547 3389
rect 1489 3380 1501 3383
rect 716 3352 1501 3380
rect 716 3340 722 3352
rect 1489 3349 1501 3352
rect 1535 3349 1547 3383
rect 2958 3380 2964 3392
rect 2919 3352 2964 3380
rect 1489 3343 1547 3349
rect 2958 3340 2964 3352
rect 3016 3340 3022 3392
rect 3786 3380 3792 3392
rect 3747 3352 3792 3380
rect 3786 3340 3792 3352
rect 3844 3340 3850 3392
rect 4154 3380 4160 3392
rect 4067 3352 4160 3380
rect 4154 3340 4160 3352
rect 4212 3380 4218 3392
rect 11698 3380 11704 3392
rect 4212 3352 11704 3380
rect 4212 3340 4218 3352
rect 11698 3340 11704 3352
rect 11756 3340 11762 3392
rect 16853 3383 16911 3389
rect 16853 3349 16865 3383
rect 16899 3380 16911 3383
rect 17494 3380 17500 3392
rect 16899 3352 17500 3380
rect 16899 3349 16911 3352
rect 16853 3343 16911 3349
rect 17494 3340 17500 3352
rect 17552 3340 17558 3392
rect 18874 3340 18880 3392
rect 18932 3380 18938 3392
rect 19337 3383 19395 3389
rect 19337 3380 19349 3383
rect 18932 3352 19349 3380
rect 18932 3340 18938 3352
rect 19337 3349 19349 3352
rect 19383 3349 19395 3383
rect 33134 3380 33140 3392
rect 33095 3352 33140 3380
rect 19337 3343 19395 3349
rect 33134 3340 33140 3352
rect 33192 3340 33198 3392
rect 1104 3290 34868 3312
rect 1104 3238 12214 3290
rect 12266 3238 12278 3290
rect 12330 3238 12342 3290
rect 12394 3238 12406 3290
rect 12458 3238 12470 3290
rect 12522 3238 23478 3290
rect 23530 3238 23542 3290
rect 23594 3238 23606 3290
rect 23658 3238 23670 3290
rect 23722 3238 23734 3290
rect 23786 3238 34868 3290
rect 1104 3216 34868 3238
rect 8021 3179 8079 3185
rect 8021 3145 8033 3179
rect 8067 3145 8079 3179
rect 13630 3176 13636 3188
rect 13591 3148 13636 3176
rect 8021 3139 8079 3145
rect 4430 3108 4436 3120
rect 1964 3080 4436 3108
rect 1964 3049 1992 3080
rect 4430 3068 4436 3080
rect 4488 3068 4494 3120
rect 1949 3043 2007 3049
rect 1949 3009 1961 3043
rect 1995 3009 2007 3043
rect 1949 3003 2007 3009
rect 2406 3000 2412 3052
rect 2464 3040 2470 3052
rect 2501 3043 2559 3049
rect 2501 3040 2513 3043
rect 2464 3012 2513 3040
rect 2464 3000 2470 3012
rect 2501 3009 2513 3012
rect 2547 3009 2559 3043
rect 4246 3040 4252 3052
rect 4207 3012 4252 3040
rect 2501 3003 2559 3009
rect 4246 3000 4252 3012
rect 4304 3000 4310 3052
rect 6822 3040 6828 3052
rect 6783 3012 6828 3040
rect 6822 3000 6828 3012
rect 6880 3000 6886 3052
rect 7742 3000 7748 3052
rect 7800 3040 7806 3052
rect 7837 3043 7895 3049
rect 7837 3040 7849 3043
rect 7800 3012 7849 3040
rect 7800 3000 7806 3012
rect 7837 3009 7849 3012
rect 7883 3009 7895 3043
rect 8036 3040 8064 3139
rect 13630 3136 13636 3148
rect 13688 3136 13694 3188
rect 13722 3136 13728 3188
rect 13780 3176 13786 3188
rect 18969 3179 19027 3185
rect 18969 3176 18981 3179
rect 13780 3148 18981 3176
rect 13780 3136 13786 3148
rect 18969 3145 18981 3148
rect 19015 3145 19027 3179
rect 19702 3176 19708 3188
rect 18969 3139 19027 3145
rect 19076 3148 19708 3176
rect 17770 3068 17776 3120
rect 17828 3108 17834 3120
rect 17865 3111 17923 3117
rect 17865 3108 17877 3111
rect 17828 3080 17877 3108
rect 17828 3068 17834 3080
rect 17865 3077 17877 3080
rect 17911 3077 17923 3111
rect 17865 3071 17923 3077
rect 18693 3111 18751 3117
rect 18693 3077 18705 3111
rect 18739 3108 18751 3111
rect 19076 3108 19104 3148
rect 19702 3136 19708 3148
rect 19760 3136 19766 3188
rect 20346 3136 20352 3188
rect 20404 3176 20410 3188
rect 22005 3179 22063 3185
rect 22005 3176 22017 3179
rect 20404 3148 22017 3176
rect 20404 3136 20410 3148
rect 22005 3145 22017 3148
rect 22051 3145 22063 3179
rect 22830 3176 22836 3188
rect 22791 3148 22836 3176
rect 22005 3139 22063 3145
rect 22830 3136 22836 3148
rect 22888 3136 22894 3188
rect 25130 3176 25136 3188
rect 25091 3148 25136 3176
rect 25130 3136 25136 3148
rect 25188 3136 25194 3188
rect 29730 3176 29736 3188
rect 29691 3148 29736 3176
rect 29730 3136 29736 3148
rect 29788 3136 29794 3188
rect 28626 3108 28632 3120
rect 18739 3080 19104 3108
rect 19168 3080 28632 3108
rect 18739 3077 18751 3080
rect 18693 3071 18751 3077
rect 8665 3043 8723 3049
rect 8665 3040 8677 3043
rect 8036 3012 8677 3040
rect 7837 3003 7895 3009
rect 8665 3009 8677 3012
rect 8711 3009 8723 3043
rect 11606 3040 11612 3052
rect 11567 3012 11612 3040
rect 8665 3003 8723 3009
rect 2225 2975 2283 2981
rect 2225 2941 2237 2975
rect 2271 2972 2283 2975
rect 2958 2972 2964 2984
rect 2271 2944 2964 2972
rect 2271 2941 2283 2944
rect 2225 2935 2283 2941
rect 2958 2932 2964 2944
rect 3016 2932 3022 2984
rect 7852 2972 7880 3003
rect 11606 3000 11612 3012
rect 11664 3000 11670 3052
rect 13538 3000 13544 3052
rect 13596 3040 13602 3052
rect 13817 3043 13875 3049
rect 13817 3040 13829 3043
rect 13596 3012 13829 3040
rect 13596 3000 13602 3012
rect 13817 3009 13829 3012
rect 13863 3009 13875 3043
rect 14366 3040 14372 3052
rect 14327 3012 14372 3040
rect 13817 3003 13875 3009
rect 14366 3000 14372 3012
rect 14424 3000 14430 3052
rect 17126 3040 17132 3052
rect 17087 3012 17132 3040
rect 17126 3000 17132 3012
rect 17184 3000 17190 3052
rect 17402 3040 17408 3052
rect 17363 3012 17408 3040
rect 17402 3000 17408 3012
rect 17460 3000 17466 3052
rect 18049 3043 18107 3049
rect 18049 3009 18061 3043
rect 18095 3040 18107 3043
rect 18322 3040 18328 3052
rect 18095 3012 18328 3040
rect 18095 3009 18107 3012
rect 18049 3003 18107 3009
rect 18322 3000 18328 3012
rect 18380 3000 18386 3052
rect 18506 3040 18512 3052
rect 18467 3012 18512 3040
rect 18506 3000 18512 3012
rect 18564 3000 18570 3052
rect 19168 3049 19196 3080
rect 28626 3068 28632 3080
rect 28684 3068 28690 3120
rect 30374 3068 30380 3120
rect 30432 3108 30438 3120
rect 30432 3080 33824 3108
rect 30432 3068 30438 3080
rect 19153 3043 19211 3049
rect 19153 3009 19165 3043
rect 19199 3009 19211 3043
rect 19153 3003 19211 3009
rect 19705 3043 19763 3049
rect 19705 3009 19717 3043
rect 19751 3040 19763 3043
rect 20165 3043 20223 3049
rect 19751 3012 20024 3040
rect 19751 3009 19763 3012
rect 19705 3003 19763 3009
rect 8297 2975 8355 2981
rect 8297 2972 8309 2975
rect 7852 2944 8309 2972
rect 8297 2941 8309 2944
rect 8343 2941 8355 2975
rect 8297 2935 8355 2941
rect 11698 2932 11704 2984
rect 11756 2972 11762 2984
rect 19242 2972 19248 2984
rect 11756 2944 19248 2972
rect 11756 2932 11762 2944
rect 19242 2932 19248 2944
rect 19300 2932 19306 2984
rect 2590 2864 2596 2916
rect 2648 2904 2654 2916
rect 3053 2907 3111 2913
rect 3053 2904 3065 2907
rect 2648 2876 3065 2904
rect 2648 2864 2654 2876
rect 3053 2873 3065 2876
rect 3099 2873 3111 2907
rect 3053 2867 3111 2873
rect 8849 2907 8907 2913
rect 8849 2873 8861 2907
rect 8895 2904 8907 2907
rect 10226 2904 10232 2916
rect 8895 2876 10232 2904
rect 8895 2873 8907 2876
rect 8849 2867 8907 2873
rect 10226 2864 10232 2876
rect 10284 2864 10290 2916
rect 10962 2864 10968 2916
rect 11020 2904 11026 2916
rect 12069 2907 12127 2913
rect 12069 2904 12081 2907
rect 11020 2876 12081 2904
rect 11020 2864 11026 2876
rect 12069 2873 12081 2876
rect 12115 2873 12127 2907
rect 12069 2867 12127 2873
rect 12434 2864 12440 2916
rect 12492 2904 12498 2916
rect 19996 2913 20024 3012
rect 20165 3009 20177 3043
rect 20211 3040 20223 3043
rect 21818 3040 21824 3052
rect 20211 3012 21824 3040
rect 20211 3009 20223 3012
rect 20165 3003 20223 3009
rect 21818 3000 21824 3012
rect 21876 3000 21882 3052
rect 21910 3000 21916 3052
rect 21968 3040 21974 3052
rect 22189 3043 22247 3049
rect 22189 3040 22201 3043
rect 21968 3012 22201 3040
rect 21968 3000 21974 3012
rect 22189 3009 22201 3012
rect 22235 3040 22247 3043
rect 22465 3043 22523 3049
rect 22465 3040 22477 3043
rect 22235 3012 22477 3040
rect 22235 3009 22247 3012
rect 22189 3003 22247 3009
rect 22465 3009 22477 3012
rect 22511 3009 22523 3043
rect 22465 3003 22523 3009
rect 24857 3043 24915 3049
rect 24857 3009 24869 3043
rect 24903 3040 24915 3043
rect 25130 3040 25136 3052
rect 24903 3012 25136 3040
rect 24903 3009 24915 3012
rect 24857 3003 24915 3009
rect 25130 3000 25136 3012
rect 25188 3000 25194 3052
rect 25498 3000 25504 3052
rect 25556 3040 25562 3052
rect 27433 3043 27491 3049
rect 27433 3040 27445 3043
rect 25556 3012 27445 3040
rect 25556 3000 25562 3012
rect 27433 3009 27445 3012
rect 27479 3040 27491 3043
rect 27709 3043 27767 3049
rect 27709 3040 27721 3043
rect 27479 3012 27721 3040
rect 27479 3009 27491 3012
rect 27433 3003 27491 3009
rect 27709 3009 27721 3012
rect 27755 3009 27767 3043
rect 27709 3003 27767 3009
rect 29638 3000 29644 3052
rect 29696 3040 29702 3052
rect 29917 3043 29975 3049
rect 29917 3040 29929 3043
rect 29696 3012 29929 3040
rect 29696 3000 29702 3012
rect 29917 3009 29929 3012
rect 29963 3040 29975 3043
rect 30193 3043 30251 3049
rect 30193 3040 30205 3043
rect 29963 3012 30205 3040
rect 29963 3009 29975 3012
rect 29917 3003 29975 3009
rect 30193 3009 30205 3012
rect 30239 3009 30251 3043
rect 30193 3003 30251 3009
rect 31294 3000 31300 3052
rect 31352 3040 31358 3052
rect 32309 3043 32367 3049
rect 32309 3040 32321 3043
rect 31352 3012 32321 3040
rect 31352 3000 31358 3012
rect 32309 3009 32321 3012
rect 32355 3009 32367 3043
rect 32309 3003 32367 3009
rect 32398 3000 32404 3052
rect 32456 3040 32462 3052
rect 33796 3049 33824 3080
rect 32953 3043 33011 3049
rect 32953 3040 32965 3043
rect 32456 3012 32965 3040
rect 32456 3000 32462 3012
rect 32953 3009 32965 3012
rect 32999 3009 33011 3043
rect 32953 3003 33011 3009
rect 33781 3043 33839 3049
rect 33781 3009 33793 3043
rect 33827 3009 33839 3043
rect 33781 3003 33839 3009
rect 28074 2972 28080 2984
rect 20732 2944 28080 2972
rect 14185 2907 14243 2913
rect 14185 2904 14197 2907
rect 12492 2876 14197 2904
rect 12492 2864 12498 2876
rect 14185 2873 14197 2876
rect 14231 2873 14243 2907
rect 14185 2867 14243 2873
rect 17589 2907 17647 2913
rect 17589 2873 17601 2907
rect 17635 2904 17647 2907
rect 19981 2907 20039 2913
rect 17635 2876 19932 2904
rect 17635 2873 17647 2876
rect 17589 2867 17647 2873
rect 1946 2796 1952 2848
rect 2004 2836 2010 2848
rect 2685 2839 2743 2845
rect 2685 2836 2697 2839
rect 2004 2808 2697 2836
rect 2004 2796 2010 2808
rect 2685 2805 2697 2808
rect 2731 2805 2743 2839
rect 2685 2799 2743 2805
rect 2866 2796 2872 2848
rect 2924 2836 2930 2848
rect 3421 2839 3479 2845
rect 3421 2836 3433 2839
rect 2924 2808 3433 2836
rect 2924 2796 2930 2808
rect 3421 2805 3433 2808
rect 3467 2805 3479 2839
rect 3421 2799 3479 2805
rect 3878 2796 3884 2848
rect 3936 2836 3942 2848
rect 4065 2839 4123 2845
rect 4065 2836 4077 2839
rect 3936 2808 4077 2836
rect 3936 2796 3942 2808
rect 4065 2805 4077 2808
rect 4111 2805 4123 2839
rect 4065 2799 4123 2805
rect 4522 2796 4528 2848
rect 4580 2836 4586 2848
rect 4709 2839 4767 2845
rect 4709 2836 4721 2839
rect 4580 2808 4721 2836
rect 4580 2796 4586 2808
rect 4709 2805 4721 2808
rect 4755 2805 4767 2839
rect 4709 2799 4767 2805
rect 5810 2796 5816 2848
rect 5868 2836 5874 2848
rect 5905 2839 5963 2845
rect 5905 2836 5917 2839
rect 5868 2808 5917 2836
rect 5868 2796 5874 2808
rect 5905 2805 5917 2808
rect 5951 2805 5963 2839
rect 5905 2799 5963 2805
rect 6454 2796 6460 2848
rect 6512 2836 6518 2848
rect 6641 2839 6699 2845
rect 6641 2836 6653 2839
rect 6512 2808 6653 2836
rect 6512 2796 6518 2808
rect 6641 2805 6653 2808
rect 6687 2805 6699 2839
rect 6641 2799 6699 2805
rect 9030 2796 9036 2848
rect 9088 2836 9094 2848
rect 9125 2839 9183 2845
rect 9125 2836 9137 2839
rect 9088 2808 9137 2836
rect 9088 2796 9094 2808
rect 9125 2805 9137 2808
rect 9171 2805 9183 2839
rect 9125 2799 9183 2805
rect 11793 2839 11851 2845
rect 11793 2805 11805 2839
rect 11839 2836 11851 2839
rect 12986 2836 12992 2848
rect 11839 2808 12992 2836
rect 11839 2805 11851 2808
rect 11793 2799 11851 2805
rect 12986 2796 12992 2808
rect 13044 2796 13050 2848
rect 13357 2839 13415 2845
rect 13357 2805 13369 2839
rect 13403 2836 13415 2839
rect 13538 2836 13544 2848
rect 13403 2808 13544 2836
rect 13403 2805 13415 2808
rect 13357 2799 13415 2805
rect 13538 2796 13544 2808
rect 13596 2796 13602 2848
rect 13722 2796 13728 2848
rect 13780 2836 13786 2848
rect 14645 2839 14703 2845
rect 14645 2836 14657 2839
rect 13780 2808 14657 2836
rect 13780 2796 13786 2808
rect 14645 2805 14657 2808
rect 14691 2805 14703 2839
rect 14645 2799 14703 2805
rect 15194 2796 15200 2848
rect 15252 2836 15258 2848
rect 16945 2839 17003 2845
rect 16945 2836 16957 2839
rect 15252 2808 16957 2836
rect 15252 2796 15258 2808
rect 16945 2805 16957 2808
rect 16991 2805 17003 2839
rect 16945 2799 17003 2805
rect 19334 2796 19340 2848
rect 19392 2836 19398 2848
rect 19521 2839 19579 2845
rect 19521 2836 19533 2839
rect 19392 2808 19533 2836
rect 19392 2796 19398 2808
rect 19521 2805 19533 2808
rect 19567 2805 19579 2839
rect 19904 2836 19932 2876
rect 19981 2873 19993 2907
rect 20027 2873 20039 2907
rect 19981 2867 20039 2873
rect 20732 2836 20760 2944
rect 28074 2932 28080 2944
rect 28132 2932 28138 2984
rect 31757 2975 31815 2981
rect 31757 2941 31769 2975
rect 31803 2972 31815 2975
rect 33502 2972 33508 2984
rect 31803 2944 33508 2972
rect 31803 2941 31815 2944
rect 31757 2935 31815 2941
rect 33502 2932 33508 2944
rect 33560 2932 33566 2984
rect 20806 2864 20812 2916
rect 20864 2904 20870 2916
rect 31297 2907 31355 2913
rect 31297 2904 31309 2907
rect 20864 2876 31309 2904
rect 20864 2864 20870 2876
rect 31297 2873 31309 2876
rect 31343 2904 31355 2907
rect 32398 2904 32404 2916
rect 31343 2876 32404 2904
rect 31343 2873 31355 2876
rect 31297 2867 31355 2873
rect 32398 2864 32404 2876
rect 32456 2864 32462 2916
rect 19904 2808 20760 2836
rect 19521 2799 19579 2805
rect 24486 2796 24492 2848
rect 24544 2836 24550 2848
rect 24673 2839 24731 2845
rect 24673 2836 24685 2839
rect 24544 2808 24685 2836
rect 24544 2796 24550 2808
rect 24673 2805 24685 2808
rect 24719 2805 24731 2839
rect 24673 2799 24731 2805
rect 27062 2796 27068 2848
rect 27120 2836 27126 2848
rect 27249 2839 27307 2845
rect 27249 2836 27261 2839
rect 27120 2808 27261 2836
rect 27120 2796 27126 2808
rect 27249 2805 27261 2808
rect 27295 2805 27307 2839
rect 29454 2836 29460 2848
rect 29415 2808 29460 2836
rect 27249 2799 27307 2805
rect 29454 2796 29460 2808
rect 29512 2796 29518 2848
rect 32214 2796 32220 2848
rect 32272 2836 32278 2848
rect 32493 2839 32551 2845
rect 32493 2836 32505 2839
rect 32272 2808 32505 2836
rect 32272 2796 32278 2808
rect 32493 2805 32505 2808
rect 32539 2805 32551 2839
rect 32493 2799 32551 2805
rect 32858 2796 32864 2848
rect 32916 2836 32922 2848
rect 33137 2839 33195 2845
rect 33137 2836 33149 2839
rect 32916 2808 33149 2836
rect 32916 2796 32922 2808
rect 33137 2805 33149 2808
rect 33183 2805 33195 2839
rect 33137 2799 33195 2805
rect 1104 2746 34868 2768
rect 1104 2694 6582 2746
rect 6634 2694 6646 2746
rect 6698 2694 6710 2746
rect 6762 2694 6774 2746
rect 6826 2694 6838 2746
rect 6890 2694 17846 2746
rect 17898 2694 17910 2746
rect 17962 2694 17974 2746
rect 18026 2694 18038 2746
rect 18090 2694 18102 2746
rect 18154 2694 29110 2746
rect 29162 2694 29174 2746
rect 29226 2694 29238 2746
rect 29290 2694 29302 2746
rect 29354 2694 29366 2746
rect 29418 2694 34868 2746
rect 1104 2672 34868 2694
rect 14366 2592 14372 2644
rect 14424 2632 14430 2644
rect 14921 2635 14979 2641
rect 14921 2632 14933 2635
rect 14424 2604 14933 2632
rect 14424 2592 14430 2604
rect 14921 2601 14933 2604
rect 14967 2601 14979 2635
rect 14921 2595 14979 2601
rect 16301 2635 16359 2641
rect 16301 2601 16313 2635
rect 16347 2632 16359 2635
rect 17310 2632 17316 2644
rect 16347 2604 17316 2632
rect 16347 2601 16359 2604
rect 16301 2595 16359 2601
rect 17310 2592 17316 2604
rect 17368 2592 17374 2644
rect 18322 2592 18328 2644
rect 18380 2632 18386 2644
rect 18380 2604 21772 2632
rect 18380 2592 18386 2604
rect 4154 2564 4160 2576
rect 3344 2536 4160 2564
rect 1394 2456 1400 2508
rect 1452 2496 1458 2508
rect 2225 2499 2283 2505
rect 2225 2496 2237 2499
rect 1452 2468 2237 2496
rect 1452 2456 1458 2468
rect 2225 2465 2237 2468
rect 2271 2496 2283 2499
rect 2590 2496 2596 2508
rect 2271 2468 2596 2496
rect 2271 2465 2283 2468
rect 2225 2459 2283 2465
rect 2590 2456 2596 2468
rect 2648 2456 2654 2508
rect 1949 2431 2007 2437
rect 1949 2397 1961 2431
rect 1995 2428 2007 2431
rect 2498 2428 2504 2440
rect 1995 2400 2504 2428
rect 1995 2397 2007 2400
rect 1949 2391 2007 2397
rect 2498 2388 2504 2400
rect 2556 2388 2562 2440
rect 2777 2431 2835 2437
rect 2777 2397 2789 2431
rect 2823 2428 2835 2431
rect 3234 2428 3240 2440
rect 2823 2400 3240 2428
rect 2823 2397 2835 2400
rect 2777 2391 2835 2397
rect 3234 2388 3240 2400
rect 3292 2388 3298 2440
rect 3344 2437 3372 2536
rect 4154 2524 4160 2536
rect 4212 2524 4218 2576
rect 6362 2524 6368 2576
rect 6420 2524 6426 2576
rect 14550 2564 14556 2576
rect 12636 2536 14556 2564
rect 3602 2456 3608 2508
rect 3660 2496 3666 2508
rect 5169 2499 5227 2505
rect 5169 2496 5181 2499
rect 3660 2468 5181 2496
rect 3660 2456 3666 2468
rect 5169 2465 5181 2468
rect 5215 2465 5227 2499
rect 6380 2496 6408 2524
rect 6641 2499 6699 2505
rect 6641 2496 6653 2499
rect 6380 2468 6653 2496
rect 5169 2459 5227 2465
rect 6641 2465 6653 2468
rect 6687 2465 6699 2499
rect 6641 2459 6699 2465
rect 7282 2456 7288 2508
rect 7340 2496 7346 2508
rect 9401 2499 9459 2505
rect 9401 2496 9413 2499
rect 7340 2468 9413 2496
rect 7340 2456 7346 2468
rect 9401 2465 9413 2468
rect 9447 2465 9459 2499
rect 9401 2459 9459 2465
rect 3329 2431 3387 2437
rect 3329 2397 3341 2431
rect 3375 2397 3387 2431
rect 3329 2391 3387 2397
rect 3418 2388 3424 2440
rect 3476 2428 3482 2440
rect 3786 2428 3792 2440
rect 3476 2400 3792 2428
rect 3476 2388 3482 2400
rect 3786 2388 3792 2400
rect 3844 2388 3850 2440
rect 4065 2431 4123 2437
rect 4065 2397 4077 2431
rect 4111 2397 4123 2431
rect 4065 2391 4123 2397
rect 2593 2363 2651 2369
rect 2593 2329 2605 2363
rect 2639 2360 2651 2363
rect 2866 2360 2872 2372
rect 2639 2332 2872 2360
rect 2639 2329 2651 2332
rect 2593 2323 2651 2329
rect 2866 2320 2872 2332
rect 2924 2320 2930 2372
rect 4080 2360 4108 2391
rect 4522 2388 4528 2440
rect 4580 2428 4586 2440
rect 4893 2431 4951 2437
rect 4893 2428 4905 2431
rect 4580 2400 4905 2428
rect 4580 2388 4586 2400
rect 4893 2397 4905 2400
rect 4939 2397 4951 2431
rect 4893 2391 4951 2397
rect 5810 2388 5816 2440
rect 5868 2428 5874 2440
rect 6365 2431 6423 2437
rect 6365 2428 6377 2431
rect 5868 2400 6377 2428
rect 5868 2388 5874 2400
rect 6365 2397 6377 2400
rect 6411 2397 6423 2431
rect 6365 2391 6423 2397
rect 7745 2431 7803 2437
rect 7745 2397 7757 2431
rect 7791 2428 7803 2431
rect 8018 2428 8024 2440
rect 7791 2400 8024 2428
rect 7791 2397 7803 2400
rect 7745 2391 7803 2397
rect 8018 2388 8024 2400
rect 8076 2388 8082 2440
rect 8110 2388 8116 2440
rect 8168 2428 8174 2440
rect 8297 2431 8355 2437
rect 8297 2428 8309 2431
rect 8168 2400 8309 2428
rect 8168 2388 8174 2400
rect 8297 2397 8309 2400
rect 8343 2397 8355 2431
rect 8297 2391 8355 2397
rect 9030 2388 9036 2440
rect 9088 2428 9094 2440
rect 9125 2431 9183 2437
rect 9125 2428 9137 2431
rect 9088 2400 9137 2428
rect 9088 2388 9094 2400
rect 9125 2397 9137 2400
rect 9171 2397 9183 2431
rect 10226 2428 10232 2440
rect 10187 2400 10232 2428
rect 9125 2391 9183 2397
rect 10226 2388 10232 2400
rect 10284 2388 10290 2440
rect 10962 2428 10968 2440
rect 10923 2400 10968 2428
rect 10962 2388 10968 2400
rect 11020 2388 11026 2440
rect 11977 2431 12035 2437
rect 11977 2397 11989 2431
rect 12023 2428 12035 2431
rect 12434 2428 12440 2440
rect 12023 2400 12440 2428
rect 12023 2397 12035 2400
rect 11977 2391 12035 2397
rect 12434 2388 12440 2400
rect 12492 2388 12498 2440
rect 12636 2437 12664 2536
rect 14550 2524 14556 2536
rect 14608 2524 14614 2576
rect 19426 2564 19432 2576
rect 18616 2536 19432 2564
rect 12986 2456 12992 2508
rect 13044 2496 13050 2508
rect 18616 2505 18644 2536
rect 19426 2524 19432 2536
rect 19484 2524 19490 2576
rect 21744 2564 21772 2604
rect 21818 2592 21824 2644
rect 21876 2632 21882 2644
rect 23293 2635 23351 2641
rect 23293 2632 23305 2635
rect 21876 2604 23305 2632
rect 21876 2592 21882 2604
rect 23293 2601 23305 2604
rect 23339 2601 23351 2635
rect 28626 2632 28632 2644
rect 28587 2604 28632 2632
rect 23293 2595 23351 2601
rect 28626 2592 28632 2604
rect 28684 2592 28690 2644
rect 31573 2567 31631 2573
rect 31573 2564 31585 2567
rect 21744 2536 31585 2564
rect 31573 2533 31585 2536
rect 31619 2533 31631 2567
rect 32950 2564 32956 2576
rect 32911 2536 32956 2564
rect 31573 2527 31631 2533
rect 32950 2524 32956 2536
rect 33008 2524 33014 2576
rect 18601 2499 18659 2505
rect 13044 2468 14320 2496
rect 13044 2456 13050 2468
rect 12621 2431 12679 2437
rect 12621 2397 12633 2431
rect 12667 2397 12679 2431
rect 12621 2391 12679 2397
rect 13449 2431 13507 2437
rect 13449 2397 13461 2431
rect 13495 2397 13507 2431
rect 13722 2428 13728 2440
rect 13683 2400 13728 2428
rect 13449 2391 13507 2397
rect 11882 2360 11888 2372
rect 4080 2332 11888 2360
rect 11882 2320 11888 2332
rect 11940 2320 11946 2372
rect 13464 2360 13492 2391
rect 13722 2388 13728 2400
rect 13780 2388 13786 2440
rect 14292 2437 14320 2468
rect 18601 2465 18613 2499
rect 18647 2465 18659 2499
rect 18601 2459 18659 2465
rect 18690 2456 18696 2508
rect 18748 2496 18754 2508
rect 19150 2496 19156 2508
rect 18748 2468 19156 2496
rect 18748 2456 18754 2468
rect 19150 2456 19156 2468
rect 19208 2496 19214 2508
rect 19245 2499 19303 2505
rect 19245 2496 19257 2499
rect 19208 2468 19257 2496
rect 19208 2456 19214 2468
rect 19245 2465 19257 2468
rect 19291 2465 19303 2499
rect 19518 2496 19524 2508
rect 19479 2468 19524 2496
rect 19245 2459 19303 2465
rect 19518 2456 19524 2468
rect 19576 2456 19582 2508
rect 20530 2456 20536 2508
rect 20588 2496 20594 2508
rect 27246 2496 27252 2508
rect 20588 2468 24440 2496
rect 27207 2468 27252 2496
rect 20588 2456 20594 2468
rect 14277 2431 14335 2437
rect 14277 2397 14289 2431
rect 14323 2397 14335 2431
rect 14277 2391 14335 2397
rect 14826 2388 14832 2440
rect 14884 2428 14890 2440
rect 15105 2431 15163 2437
rect 15105 2428 15117 2431
rect 14884 2400 15117 2428
rect 14884 2388 14890 2400
rect 15105 2397 15117 2400
rect 15151 2428 15163 2431
rect 15381 2431 15439 2437
rect 15381 2428 15393 2431
rect 15151 2400 15393 2428
rect 15151 2397 15163 2400
rect 15105 2391 15163 2397
rect 15381 2397 15393 2400
rect 15427 2397 15439 2431
rect 15381 2391 15439 2397
rect 15841 2431 15899 2437
rect 15841 2397 15853 2431
rect 15887 2428 15899 2431
rect 16117 2431 16175 2437
rect 16117 2428 16129 2431
rect 15887 2400 16129 2428
rect 15887 2397 15899 2400
rect 15841 2391 15899 2397
rect 16117 2397 16129 2400
rect 16163 2428 16175 2431
rect 16758 2428 16764 2440
rect 16163 2400 16764 2428
rect 16163 2397 16175 2400
rect 16117 2391 16175 2397
rect 16758 2388 16764 2400
rect 16816 2388 16822 2440
rect 16942 2428 16948 2440
rect 16903 2400 16948 2428
rect 16942 2388 16948 2400
rect 17000 2388 17006 2440
rect 17494 2428 17500 2440
rect 17455 2400 17500 2428
rect 17494 2388 17500 2400
rect 17552 2388 17558 2440
rect 18046 2388 18052 2440
rect 18104 2428 18110 2440
rect 18874 2428 18880 2440
rect 18104 2400 18880 2428
rect 18104 2388 18110 2400
rect 18874 2388 18880 2400
rect 18932 2388 18938 2440
rect 20625 2431 20683 2437
rect 20625 2397 20637 2431
rect 20671 2428 20683 2431
rect 20901 2431 20959 2437
rect 20901 2428 20913 2431
rect 20671 2400 20913 2428
rect 20671 2397 20683 2400
rect 20625 2391 20683 2397
rect 20901 2397 20913 2400
rect 20947 2397 20959 2431
rect 22094 2428 22100 2440
rect 22055 2400 22100 2428
rect 20901 2391 20959 2397
rect 16850 2360 16856 2372
rect 13464 2332 16856 2360
rect 16850 2320 16856 2332
rect 16908 2320 16914 2372
rect 18782 2320 18788 2372
rect 18840 2360 18846 2372
rect 20640 2360 20668 2391
rect 22094 2388 22100 2400
rect 22152 2388 22158 2440
rect 22830 2388 22836 2440
rect 22888 2428 22894 2440
rect 22925 2431 22983 2437
rect 22925 2428 22937 2431
rect 22888 2400 22937 2428
rect 22888 2388 22894 2400
rect 22925 2397 22937 2400
rect 22971 2397 22983 2431
rect 23474 2428 23480 2440
rect 23435 2400 23480 2428
rect 22925 2391 22983 2397
rect 23474 2388 23480 2400
rect 23532 2428 23538 2440
rect 24412 2437 24440 2468
rect 27246 2456 27252 2468
rect 27304 2456 27310 2508
rect 29822 2496 29828 2508
rect 29783 2468 29828 2496
rect 29822 2456 29828 2468
rect 29880 2456 29886 2508
rect 31846 2456 31852 2508
rect 31904 2496 31910 2508
rect 33505 2499 33563 2505
rect 31904 2468 32536 2496
rect 31904 2456 31910 2468
rect 23753 2431 23811 2437
rect 23753 2428 23765 2431
rect 23532 2400 23765 2428
rect 23532 2388 23538 2400
rect 23753 2397 23765 2400
rect 23799 2397 23811 2431
rect 23753 2391 23811 2397
rect 24397 2431 24455 2437
rect 24397 2397 24409 2431
rect 24443 2397 24455 2431
rect 25222 2428 25228 2440
rect 25183 2400 25228 2428
rect 24397 2391 24455 2397
rect 25222 2388 25228 2400
rect 25280 2388 25286 2440
rect 26973 2431 27031 2437
rect 26973 2428 26985 2431
rect 26528 2400 26985 2428
rect 18840 2332 20668 2360
rect 18840 2320 18846 2332
rect 2774 2252 2780 2304
rect 2832 2292 2838 2304
rect 3145 2295 3203 2301
rect 3145 2292 3157 2295
rect 2832 2264 3157 2292
rect 2832 2252 2838 2264
rect 3145 2261 3157 2264
rect 3191 2261 3203 2295
rect 3145 2255 3203 2261
rect 7098 2252 7104 2304
rect 7156 2292 7162 2304
rect 7561 2295 7619 2301
rect 7561 2292 7573 2295
rect 7156 2264 7573 2292
rect 7156 2252 7162 2264
rect 7561 2261 7573 2264
rect 7607 2261 7619 2295
rect 7561 2255 7619 2261
rect 8386 2252 8392 2304
rect 8444 2292 8450 2304
rect 8481 2295 8539 2301
rect 8481 2292 8493 2295
rect 8444 2264 8493 2292
rect 8444 2252 8450 2264
rect 8481 2261 8493 2264
rect 8527 2261 8539 2295
rect 8481 2255 8539 2261
rect 9674 2252 9680 2304
rect 9732 2292 9738 2304
rect 10413 2295 10471 2301
rect 10413 2292 10425 2295
rect 9732 2264 10425 2292
rect 9732 2252 9738 2264
rect 10413 2261 10425 2264
rect 10459 2261 10471 2295
rect 11146 2292 11152 2304
rect 11107 2264 11152 2292
rect 10413 2255 10471 2261
rect 11146 2252 11152 2264
rect 11204 2252 11210 2304
rect 11606 2252 11612 2304
rect 11664 2292 11670 2304
rect 11793 2295 11851 2301
rect 11793 2292 11805 2295
rect 11664 2264 11805 2292
rect 11664 2252 11670 2264
rect 11793 2261 11805 2264
rect 11839 2261 11851 2295
rect 11793 2255 11851 2261
rect 12066 2252 12072 2304
rect 12124 2292 12130 2304
rect 12437 2295 12495 2301
rect 12437 2292 12449 2295
rect 12124 2264 12449 2292
rect 12124 2252 12130 2264
rect 12437 2261 12449 2264
rect 12483 2261 12495 2295
rect 12437 2255 12495 2261
rect 12894 2252 12900 2304
rect 12952 2292 12958 2304
rect 13722 2292 13728 2304
rect 12952 2264 13728 2292
rect 12952 2252 12958 2264
rect 13722 2252 13728 2264
rect 13780 2252 13786 2304
rect 14182 2252 14188 2304
rect 14240 2292 14246 2304
rect 14461 2295 14519 2301
rect 14461 2292 14473 2295
rect 14240 2264 14473 2292
rect 14240 2252 14246 2264
rect 14461 2261 14473 2264
rect 14507 2261 14519 2295
rect 14461 2255 14519 2261
rect 16114 2252 16120 2304
rect 16172 2292 16178 2304
rect 16761 2295 16819 2301
rect 16761 2292 16773 2295
rect 16172 2264 16773 2292
rect 16172 2252 16178 2264
rect 16761 2261 16773 2264
rect 16807 2261 16819 2295
rect 16761 2255 16819 2261
rect 17402 2252 17408 2304
rect 17460 2292 17466 2304
rect 17681 2295 17739 2301
rect 17681 2292 17693 2295
rect 17460 2264 17693 2292
rect 17460 2252 17466 2264
rect 17681 2261 17693 2264
rect 17727 2261 17739 2295
rect 17681 2255 17739 2261
rect 19978 2252 19984 2304
rect 20036 2292 20042 2304
rect 20441 2295 20499 2301
rect 20441 2292 20453 2295
rect 20036 2264 20453 2292
rect 20036 2252 20042 2264
rect 20441 2261 20453 2264
rect 20487 2261 20499 2295
rect 20441 2255 20499 2261
rect 21266 2252 21272 2304
rect 21324 2292 21330 2304
rect 21913 2295 21971 2301
rect 21913 2292 21925 2295
rect 21324 2264 21925 2292
rect 21324 2252 21330 2264
rect 21913 2261 21925 2264
rect 21959 2261 21971 2295
rect 21913 2255 21971 2261
rect 22554 2252 22560 2304
rect 22612 2292 22618 2304
rect 22741 2295 22799 2301
rect 22741 2292 22753 2295
rect 22612 2264 22753 2292
rect 22612 2252 22618 2264
rect 22741 2261 22753 2264
rect 22787 2261 22799 2295
rect 22741 2255 22799 2261
rect 23842 2252 23848 2304
rect 23900 2292 23906 2304
rect 24581 2295 24639 2301
rect 24581 2292 24593 2295
rect 23900 2264 24593 2292
rect 23900 2252 23906 2264
rect 24581 2261 24593 2264
rect 24627 2261 24639 2295
rect 24581 2255 24639 2261
rect 25130 2252 25136 2304
rect 25188 2292 25194 2304
rect 25409 2295 25467 2301
rect 25409 2292 25421 2295
rect 25188 2264 25421 2292
rect 25188 2252 25194 2264
rect 25409 2261 25421 2264
rect 25455 2261 25467 2295
rect 25409 2255 25467 2261
rect 26418 2252 26424 2304
rect 26476 2292 26482 2304
rect 26528 2301 26556 2400
rect 26973 2397 26985 2400
rect 27019 2397 27031 2431
rect 28074 2428 28080 2440
rect 28035 2400 28080 2428
rect 26973 2391 27031 2397
rect 28074 2388 28080 2400
rect 28132 2388 28138 2440
rect 28350 2388 28356 2440
rect 28408 2428 28414 2440
rect 28813 2431 28871 2437
rect 28813 2428 28825 2431
rect 28408 2400 28825 2428
rect 28408 2388 28414 2400
rect 28813 2397 28825 2400
rect 28859 2397 28871 2431
rect 28813 2391 28871 2397
rect 28828 2360 28856 2391
rect 28994 2388 29000 2440
rect 29052 2428 29058 2440
rect 29454 2428 29460 2440
rect 29052 2400 29460 2428
rect 29052 2388 29058 2400
rect 29454 2388 29460 2400
rect 29512 2428 29518 2440
rect 29549 2431 29607 2437
rect 29549 2428 29561 2431
rect 29512 2400 29561 2428
rect 29512 2388 29518 2400
rect 29549 2397 29561 2400
rect 29595 2397 29607 2431
rect 30926 2428 30932 2440
rect 30887 2400 30932 2428
rect 29549 2391 29607 2397
rect 30926 2388 30932 2400
rect 30984 2388 30990 2440
rect 31297 2431 31355 2437
rect 31297 2397 31309 2431
rect 31343 2428 31355 2431
rect 31570 2428 31576 2440
rect 31343 2400 31576 2428
rect 31343 2397 31355 2400
rect 31297 2391 31355 2397
rect 31570 2388 31576 2400
rect 31628 2428 31634 2440
rect 31757 2431 31815 2437
rect 31757 2428 31769 2431
rect 31628 2400 31769 2428
rect 31628 2388 31634 2400
rect 31757 2397 31769 2400
rect 31803 2397 31815 2431
rect 32398 2428 32404 2440
rect 32359 2400 32404 2428
rect 31757 2391 31815 2397
rect 32398 2388 32404 2400
rect 32456 2388 32462 2440
rect 32508 2428 32536 2468
rect 33505 2465 33517 2499
rect 33551 2496 33563 2499
rect 33870 2496 33876 2508
rect 33551 2468 33876 2496
rect 33551 2465 33563 2468
rect 33505 2459 33563 2465
rect 33870 2456 33876 2468
rect 33928 2456 33934 2508
rect 33781 2431 33839 2437
rect 33781 2428 33793 2431
rect 32508 2400 33793 2428
rect 33781 2397 33793 2400
rect 33827 2397 33839 2431
rect 33781 2391 33839 2397
rect 29089 2363 29147 2369
rect 29089 2360 29101 2363
rect 28828 2332 29101 2360
rect 29089 2329 29101 2332
rect 29135 2329 29147 2363
rect 33134 2360 33140 2372
rect 33095 2332 33140 2360
rect 29089 2323 29147 2329
rect 33134 2320 33140 2332
rect 33192 2320 33198 2372
rect 26513 2295 26571 2301
rect 26513 2292 26525 2295
rect 26476 2264 26525 2292
rect 26476 2252 26482 2264
rect 26513 2261 26525 2264
rect 26559 2261 26571 2295
rect 26513 2255 26571 2261
rect 27706 2252 27712 2304
rect 27764 2292 27770 2304
rect 28261 2295 28319 2301
rect 28261 2292 28273 2295
rect 27764 2264 28273 2292
rect 27764 2252 27770 2264
rect 28261 2261 28273 2264
rect 28307 2261 28319 2295
rect 28261 2255 28319 2261
rect 30282 2252 30288 2304
rect 30340 2292 30346 2304
rect 30745 2295 30803 2301
rect 30745 2292 30757 2295
rect 30340 2264 30757 2292
rect 30340 2252 30346 2264
rect 30745 2261 30757 2264
rect 30791 2261 30803 2295
rect 32582 2292 32588 2304
rect 32543 2264 32588 2292
rect 30745 2255 30803 2261
rect 32582 2252 32588 2264
rect 32640 2252 32646 2304
rect 1104 2202 34868 2224
rect 1104 2150 12214 2202
rect 12266 2150 12278 2202
rect 12330 2150 12342 2202
rect 12394 2150 12406 2202
rect 12458 2150 12470 2202
rect 12522 2150 23478 2202
rect 23530 2150 23542 2202
rect 23594 2150 23606 2202
rect 23658 2150 23670 2202
rect 23722 2150 23734 2202
rect 23786 2150 34868 2202
rect 1104 2128 34868 2150
rect 2498 2048 2504 2100
rect 2556 2088 2562 2100
rect 2556 2060 11744 2088
rect 2556 2048 2562 2060
rect 3234 1980 3240 2032
rect 3292 2020 3298 2032
rect 11716 2020 11744 2060
rect 11882 2048 11888 2100
rect 11940 2088 11946 2100
rect 17218 2088 17224 2100
rect 11940 2060 17224 2088
rect 11940 2048 11946 2060
rect 17218 2048 17224 2060
rect 17276 2048 17282 2100
rect 16666 2020 16672 2032
rect 3292 1992 6914 2020
rect 11716 1992 16672 2020
rect 3292 1980 3298 1992
rect 6886 1884 6914 1992
rect 16666 1980 16672 1992
rect 16724 1980 16730 2032
rect 11146 1912 11152 1964
rect 11204 1952 11210 1964
rect 18506 1952 18512 1964
rect 11204 1924 18512 1952
rect 11204 1912 11210 1924
rect 18506 1912 18512 1924
rect 18564 1912 18570 1964
rect 18230 1884 18236 1896
rect 6886 1856 18236 1884
rect 18230 1844 18236 1856
rect 18288 1844 18294 1896
rect 8018 1776 8024 1828
rect 8076 1816 8082 1828
rect 15194 1816 15200 1828
rect 8076 1788 15200 1816
rect 8076 1776 8082 1788
rect 15194 1776 15200 1788
rect 15252 1776 15258 1828
<< via1 >>
rect 11612 33940 11664 33992
rect 18420 33940 18472 33992
rect 10508 33872 10560 33924
rect 15016 33872 15068 33924
rect 16672 33872 16724 33924
rect 20260 33872 20312 33924
rect 14372 33804 14424 33856
rect 18972 33804 19024 33856
rect 12214 33702 12266 33754
rect 12278 33702 12330 33754
rect 12342 33702 12394 33754
rect 12406 33702 12458 33754
rect 12470 33702 12522 33754
rect 23478 33702 23530 33754
rect 23542 33702 23594 33754
rect 23606 33702 23658 33754
rect 23670 33702 23722 33754
rect 23734 33702 23786 33754
rect 3884 33600 3936 33652
rect 6736 33643 6788 33652
rect 6736 33609 6745 33643
rect 6745 33609 6779 33643
rect 6779 33609 6788 33643
rect 6736 33600 6788 33609
rect 9864 33643 9916 33652
rect 9864 33609 9873 33643
rect 9873 33609 9907 33643
rect 9907 33609 9916 33643
rect 9864 33600 9916 33609
rect 2780 33575 2832 33584
rect 2780 33541 2789 33575
rect 2789 33541 2823 33575
rect 2823 33541 2832 33575
rect 2780 33532 2832 33541
rect 16672 33600 16724 33652
rect 16764 33600 16816 33652
rect 18052 33600 18104 33652
rect 23020 33643 23072 33652
rect 23020 33609 23029 33643
rect 23029 33609 23063 33643
rect 23063 33609 23072 33643
rect 23020 33600 23072 33609
rect 23940 33643 23992 33652
rect 23940 33609 23949 33643
rect 23949 33609 23983 33643
rect 23983 33609 23992 33643
rect 23940 33600 23992 33609
rect 26056 33643 26108 33652
rect 26056 33609 26065 33643
rect 26065 33609 26099 33643
rect 26099 33609 26108 33643
rect 26056 33600 26108 33609
rect 26516 33643 26568 33652
rect 26516 33609 26525 33643
rect 26525 33609 26559 33643
rect 26559 33609 26568 33643
rect 26516 33600 26568 33609
rect 28172 33643 28224 33652
rect 28172 33609 28181 33643
rect 28181 33609 28215 33643
rect 28215 33609 28224 33643
rect 28172 33600 28224 33609
rect 29092 33643 29144 33652
rect 29092 33609 29101 33643
rect 29101 33609 29135 33643
rect 29135 33609 29144 33643
rect 29092 33600 29144 33609
rect 29920 33643 29972 33652
rect 29920 33609 29929 33643
rect 29929 33609 29963 33643
rect 29963 33609 29972 33643
rect 29920 33600 29972 33609
rect 31760 33643 31812 33652
rect 31760 33609 31769 33643
rect 31769 33609 31803 33643
rect 31803 33609 31812 33643
rect 31760 33600 31812 33609
rect 1032 33464 1084 33516
rect 2228 33507 2280 33516
rect 2228 33473 2237 33507
rect 2237 33473 2271 33507
rect 2271 33473 2280 33507
rect 2228 33464 2280 33473
rect 3976 33507 4028 33516
rect 3976 33473 3985 33507
rect 3985 33473 4019 33507
rect 4019 33473 4028 33507
rect 4620 33507 4672 33516
rect 3976 33464 4028 33473
rect 4620 33473 4629 33507
rect 4629 33473 4663 33507
rect 4663 33473 4672 33507
rect 4620 33464 4672 33473
rect 5540 33464 5592 33516
rect 6368 33464 6420 33516
rect 7932 33507 7984 33516
rect 7932 33473 7941 33507
rect 7941 33473 7975 33507
rect 7975 33473 7984 33507
rect 7932 33464 7984 33473
rect 8484 33464 8536 33516
rect 14740 33532 14792 33584
rect 15476 33532 15528 33584
rect 11704 33507 11756 33516
rect 3056 33396 3108 33448
rect 10508 33396 10560 33448
rect 10600 33396 10652 33448
rect 11152 33439 11204 33448
rect 11152 33405 11161 33439
rect 11161 33405 11195 33439
rect 11195 33405 11204 33439
rect 11152 33396 11204 33405
rect 11704 33473 11713 33507
rect 11713 33473 11747 33507
rect 11747 33473 11756 33507
rect 11704 33464 11756 33473
rect 14372 33507 14424 33516
rect 14372 33473 14381 33507
rect 14381 33473 14415 33507
rect 14415 33473 14424 33507
rect 14372 33464 14424 33473
rect 14464 33464 14516 33516
rect 18604 33532 18656 33584
rect 17132 33507 17184 33516
rect 11612 33328 11664 33380
rect 2596 33260 2648 33312
rect 3976 33260 4028 33312
rect 8024 33303 8076 33312
rect 8024 33269 8033 33303
rect 8033 33269 8067 33303
rect 8067 33269 8076 33303
rect 8024 33260 8076 33269
rect 11888 33303 11940 33312
rect 11888 33269 11897 33303
rect 11897 33269 11931 33303
rect 11931 33269 11940 33303
rect 11888 33260 11940 33269
rect 13820 33328 13872 33380
rect 17132 33473 17141 33507
rect 17141 33473 17175 33507
rect 17175 33473 17184 33507
rect 17132 33464 17184 33473
rect 18788 33464 18840 33516
rect 19432 33507 19484 33516
rect 19432 33473 19441 33507
rect 19441 33473 19475 33507
rect 19475 33473 19484 33507
rect 19432 33464 19484 33473
rect 20628 33507 20680 33516
rect 20628 33473 20637 33507
rect 20637 33473 20671 33507
rect 20671 33473 20680 33507
rect 20628 33464 20680 33473
rect 21272 33464 21324 33516
rect 25872 33507 25924 33516
rect 25872 33473 25881 33507
rect 25881 33473 25915 33507
rect 25915 33473 25924 33507
rect 25872 33464 25924 33473
rect 28724 33464 28776 33516
rect 30380 33507 30432 33516
rect 17408 33396 17460 33448
rect 19800 33396 19852 33448
rect 24492 33396 24544 33448
rect 27344 33396 27396 33448
rect 27620 33396 27672 33448
rect 30380 33473 30389 33507
rect 30389 33473 30423 33507
rect 30423 33473 30432 33507
rect 30380 33464 30432 33473
rect 33324 33464 33376 33516
rect 34428 33464 34480 33516
rect 31208 33396 31260 33448
rect 33232 33396 33284 33448
rect 33600 33396 33652 33448
rect 33784 33439 33836 33448
rect 33784 33405 33793 33439
rect 33793 33405 33827 33439
rect 33827 33405 33836 33439
rect 33784 33396 33836 33405
rect 15568 33260 15620 33312
rect 17776 33328 17828 33380
rect 19340 33328 19392 33380
rect 32312 33371 32364 33380
rect 32312 33337 32321 33371
rect 32321 33337 32355 33371
rect 32355 33337 32364 33371
rect 32312 33328 32364 33337
rect 32864 33328 32916 33380
rect 18512 33260 18564 33312
rect 21916 33260 21968 33312
rect 30840 33260 30892 33312
rect 6582 33158 6634 33210
rect 6646 33158 6698 33210
rect 6710 33158 6762 33210
rect 6774 33158 6826 33210
rect 6838 33158 6890 33210
rect 17846 33158 17898 33210
rect 17910 33158 17962 33210
rect 17974 33158 18026 33210
rect 18038 33158 18090 33210
rect 18102 33158 18154 33210
rect 29110 33158 29162 33210
rect 29174 33158 29226 33210
rect 29238 33158 29290 33210
rect 29302 33158 29354 33210
rect 29366 33158 29418 33210
rect 2228 33056 2280 33108
rect 4620 33056 4672 33108
rect 5540 33099 5592 33108
rect 5540 33065 5549 33099
rect 5549 33065 5583 33099
rect 5583 33065 5592 33099
rect 5540 33056 5592 33065
rect 6000 33099 6052 33108
rect 6000 33065 6009 33099
rect 6009 33065 6043 33099
rect 6043 33065 6052 33099
rect 6000 33056 6052 33065
rect 8484 33099 8536 33108
rect 8484 33065 8493 33099
rect 8493 33065 8527 33099
rect 8527 33065 8536 33099
rect 8484 33056 8536 33065
rect 10784 33099 10836 33108
rect 10784 33065 10793 33099
rect 10793 33065 10827 33099
rect 10827 33065 10836 33099
rect 10784 33056 10836 33065
rect 11152 33056 11204 33108
rect 14648 33099 14700 33108
rect 14648 33065 14657 33099
rect 14657 33065 14691 33099
rect 14691 33065 14700 33099
rect 14648 33056 14700 33065
rect 16396 33099 16448 33108
rect 16396 33065 16405 33099
rect 16405 33065 16439 33099
rect 16439 33065 16448 33099
rect 16396 33056 16448 33065
rect 17132 33056 17184 33108
rect 18696 33056 18748 33108
rect 20628 33056 20680 33108
rect 24676 33099 24728 33108
rect 1308 32988 1360 33040
rect 14740 32988 14792 33040
rect 15016 32920 15068 32972
rect 20 32852 72 32904
rect 1308 32852 1360 32904
rect 2136 32852 2188 32904
rect 2780 32852 2832 32904
rect 3516 32852 3568 32904
rect 9312 32895 9364 32904
rect 1860 32827 1912 32836
rect 1860 32793 1869 32827
rect 1869 32793 1903 32827
rect 1903 32793 1912 32827
rect 1860 32784 1912 32793
rect 9312 32861 9321 32895
rect 9321 32861 9355 32895
rect 9355 32861 9364 32895
rect 9312 32852 9364 32861
rect 10784 32852 10836 32904
rect 15200 32895 15252 32904
rect 15200 32861 15209 32895
rect 15209 32861 15243 32895
rect 15243 32861 15252 32895
rect 15200 32852 15252 32861
rect 15568 32852 15620 32904
rect 24676 33065 24685 33099
rect 24685 33065 24719 33099
rect 24719 33065 24728 33099
rect 24676 33056 24728 33065
rect 25412 33099 25464 33108
rect 25412 33065 25421 33099
rect 25421 33065 25455 33099
rect 25455 33065 25464 33099
rect 25412 33056 25464 33065
rect 27252 33099 27304 33108
rect 27252 33065 27261 33099
rect 27261 33065 27295 33099
rect 27295 33065 27304 33099
rect 27252 33056 27304 33065
rect 30380 33056 30432 33108
rect 30748 33099 30800 33108
rect 30748 33065 30757 33099
rect 30757 33065 30791 33099
rect 30791 33065 30800 33099
rect 30748 33056 30800 33065
rect 32496 33099 32548 33108
rect 32496 33065 32505 33099
rect 32505 33065 32539 33099
rect 32539 33065 32548 33099
rect 32496 33056 32548 33065
rect 33140 33099 33192 33108
rect 33140 33065 33149 33099
rect 33149 33065 33183 33099
rect 33183 33065 33192 33099
rect 33140 33056 33192 33065
rect 33692 33099 33744 33108
rect 33692 33065 33701 33099
rect 33701 33065 33735 33099
rect 33735 33065 33744 33099
rect 33692 33056 33744 33065
rect 19248 32895 19300 32904
rect 15292 32784 15344 32836
rect 18512 32827 18564 32836
rect 18512 32793 18521 32827
rect 18521 32793 18555 32827
rect 18555 32793 18564 32827
rect 18512 32784 18564 32793
rect 19248 32861 19257 32895
rect 19257 32861 19291 32895
rect 19291 32861 19300 32895
rect 19248 32852 19300 32861
rect 21916 32895 21968 32904
rect 21916 32861 21925 32895
rect 21925 32861 21959 32895
rect 21959 32861 21968 32895
rect 21916 32852 21968 32861
rect 33784 32988 33836 33040
rect 19340 32784 19392 32836
rect 29920 32920 29972 32972
rect 30748 32920 30800 32972
rect 31944 32920 31996 32972
rect 27896 32895 27948 32904
rect 27896 32861 27905 32895
rect 27905 32861 27939 32895
rect 27939 32861 27948 32895
rect 31300 32895 31352 32904
rect 27896 32852 27948 32861
rect 31300 32861 31309 32895
rect 31309 32861 31343 32895
rect 31343 32861 31352 32895
rect 31300 32852 31352 32861
rect 32956 32895 33008 32904
rect 32956 32861 32965 32895
rect 32965 32861 32999 32895
rect 32999 32861 33008 32895
rect 32956 32852 33008 32861
rect 34244 32895 34296 32904
rect 34244 32861 34253 32895
rect 34253 32861 34287 32895
rect 34287 32861 34296 32895
rect 34244 32852 34296 32861
rect 2320 32759 2372 32768
rect 2320 32725 2329 32759
rect 2329 32725 2363 32759
rect 2363 32725 2372 32759
rect 2320 32716 2372 32725
rect 6460 32759 6512 32768
rect 6460 32725 6469 32759
rect 6469 32725 6503 32759
rect 6503 32725 6512 32759
rect 6460 32716 6512 32725
rect 9128 32759 9180 32768
rect 9128 32725 9137 32759
rect 9137 32725 9171 32759
rect 9171 32725 9180 32759
rect 9128 32716 9180 32725
rect 11244 32759 11296 32768
rect 11244 32725 11253 32759
rect 11253 32725 11287 32759
rect 11287 32725 11296 32759
rect 11244 32716 11296 32725
rect 32772 32784 32824 32836
rect 28724 32759 28776 32768
rect 28724 32725 28733 32759
rect 28733 32725 28767 32759
rect 28767 32725 28776 32759
rect 28724 32716 28776 32725
rect 28816 32716 28868 32768
rect 12214 32614 12266 32666
rect 12278 32614 12330 32666
rect 12342 32614 12394 32666
rect 12406 32614 12458 32666
rect 12470 32614 12522 32666
rect 23478 32614 23530 32666
rect 23542 32614 23594 32666
rect 23606 32614 23658 32666
rect 23670 32614 23722 32666
rect 23734 32614 23786 32666
rect 2872 32512 2924 32564
rect 15568 32555 15620 32564
rect 15568 32521 15577 32555
rect 15577 32521 15611 32555
rect 15611 32521 15620 32555
rect 15568 32512 15620 32521
rect 24860 32512 24912 32564
rect 28816 32512 28868 32564
rect 32772 32555 32824 32564
rect 32772 32521 32781 32555
rect 32781 32521 32815 32555
rect 32815 32521 32824 32555
rect 32772 32512 32824 32521
rect 1308 32444 1360 32496
rect 11244 32376 11296 32428
rect 18512 32419 18564 32428
rect 18512 32385 18521 32419
rect 18521 32385 18555 32419
rect 18555 32385 18564 32419
rect 18512 32376 18564 32385
rect 27896 32444 27948 32496
rect 34152 32512 34204 32564
rect 30380 32376 30432 32428
rect 33416 32376 33468 32428
rect 1400 32351 1452 32360
rect 1400 32317 1409 32351
rect 1409 32317 1443 32351
rect 1443 32317 1452 32351
rect 1400 32308 1452 32317
rect 1768 32308 1820 32360
rect 33324 32308 33376 32360
rect 33600 32376 33652 32428
rect 31944 32172 31996 32224
rect 34244 32215 34296 32224
rect 34244 32181 34253 32215
rect 34253 32181 34287 32215
rect 34287 32181 34296 32215
rect 34244 32172 34296 32181
rect 6582 32070 6634 32122
rect 6646 32070 6698 32122
rect 6710 32070 6762 32122
rect 6774 32070 6826 32122
rect 6838 32070 6890 32122
rect 17846 32070 17898 32122
rect 17910 32070 17962 32122
rect 17974 32070 18026 32122
rect 18038 32070 18090 32122
rect 18102 32070 18154 32122
rect 29110 32070 29162 32122
rect 29174 32070 29226 32122
rect 29238 32070 29290 32122
rect 29302 32070 29354 32122
rect 29366 32070 29418 32122
rect 2964 31968 3016 32020
rect 33232 31968 33284 32020
rect 33416 31968 33468 32020
rect 35440 31968 35492 32020
rect 2780 31900 2832 31952
rect 1676 31807 1728 31816
rect 1676 31773 1685 31807
rect 1685 31773 1719 31807
rect 1719 31773 1728 31807
rect 1676 31764 1728 31773
rect 2964 31807 3016 31816
rect 2964 31773 2973 31807
rect 2973 31773 3007 31807
rect 3007 31773 3016 31807
rect 2964 31764 3016 31773
rect 32956 31764 33008 31816
rect 33600 31807 33652 31816
rect 33600 31773 33609 31807
rect 33609 31773 33643 31807
rect 33643 31773 33652 31807
rect 33600 31764 33652 31773
rect 1492 31671 1544 31680
rect 1492 31637 1501 31671
rect 1501 31637 1535 31671
rect 1535 31637 1544 31671
rect 1492 31628 1544 31637
rect 12214 31526 12266 31578
rect 12278 31526 12330 31578
rect 12342 31526 12394 31578
rect 12406 31526 12458 31578
rect 12470 31526 12522 31578
rect 23478 31526 23530 31578
rect 23542 31526 23594 31578
rect 23606 31526 23658 31578
rect 23670 31526 23722 31578
rect 23734 31526 23786 31578
rect 1400 31467 1452 31476
rect 1400 31433 1409 31467
rect 1409 31433 1443 31467
rect 1443 31433 1452 31467
rect 1400 31424 1452 31433
rect 11888 31356 11940 31408
rect 34336 31331 34388 31340
rect 34336 31297 34345 31331
rect 34345 31297 34379 31331
rect 34379 31297 34388 31331
rect 34336 31288 34388 31297
rect 22100 31084 22152 31136
rect 33416 31127 33468 31136
rect 33416 31093 33425 31127
rect 33425 31093 33459 31127
rect 33459 31093 33468 31127
rect 33416 31084 33468 31093
rect 33692 31084 33744 31136
rect 6582 30982 6634 31034
rect 6646 30982 6698 31034
rect 6710 30982 6762 31034
rect 6774 30982 6826 31034
rect 6838 30982 6890 31034
rect 17846 30982 17898 31034
rect 17910 30982 17962 31034
rect 17974 30982 18026 31034
rect 18038 30982 18090 31034
rect 18102 30982 18154 31034
rect 29110 30982 29162 31034
rect 29174 30982 29226 31034
rect 29238 30982 29290 31034
rect 29302 30982 29354 31034
rect 29366 30982 29418 31034
rect 22100 30880 22152 30932
rect 34060 30880 34112 30932
rect 30380 30744 30432 30796
rect 34336 30719 34388 30728
rect 1492 30583 1544 30592
rect 1492 30549 1501 30583
rect 1501 30549 1535 30583
rect 1535 30549 1544 30583
rect 1492 30540 1544 30549
rect 34336 30685 34345 30719
rect 34345 30685 34379 30719
rect 34379 30685 34388 30719
rect 34336 30676 34388 30685
rect 2136 30540 2188 30592
rect 12214 30438 12266 30490
rect 12278 30438 12330 30490
rect 12342 30438 12394 30490
rect 12406 30438 12458 30490
rect 12470 30438 12522 30490
rect 23478 30438 23530 30490
rect 23542 30438 23594 30490
rect 23606 30438 23658 30490
rect 23670 30438 23722 30490
rect 23734 30438 23786 30490
rect 34336 30336 34388 30388
rect 34336 30243 34388 30252
rect 34336 30209 34345 30243
rect 34345 30209 34379 30243
rect 34379 30209 34388 30243
rect 34336 30200 34388 30209
rect 1952 30064 2004 30116
rect 18512 30132 18564 30184
rect 33876 29996 33928 30048
rect 6582 29894 6634 29946
rect 6646 29894 6698 29946
rect 6710 29894 6762 29946
rect 6774 29894 6826 29946
rect 6838 29894 6890 29946
rect 17846 29894 17898 29946
rect 17910 29894 17962 29946
rect 17974 29894 18026 29946
rect 18038 29894 18090 29946
rect 18102 29894 18154 29946
rect 29110 29894 29162 29946
rect 29174 29894 29226 29946
rect 29238 29894 29290 29946
rect 29302 29894 29354 29946
rect 29366 29894 29418 29946
rect 1952 29835 2004 29844
rect 1952 29801 1961 29835
rect 1961 29801 1995 29835
rect 1995 29801 2004 29835
rect 1952 29792 2004 29801
rect 33600 29792 33652 29844
rect 34336 29631 34388 29640
rect 34336 29597 34345 29631
rect 34345 29597 34379 29631
rect 34379 29597 34388 29631
rect 34336 29588 34388 29597
rect 1492 29495 1544 29504
rect 1492 29461 1501 29495
rect 1501 29461 1535 29495
rect 1535 29461 1544 29495
rect 1492 29452 1544 29461
rect 2412 29495 2464 29504
rect 2412 29461 2421 29495
rect 2421 29461 2455 29495
rect 2455 29461 2464 29495
rect 2412 29452 2464 29461
rect 12214 29350 12266 29402
rect 12278 29350 12330 29402
rect 12342 29350 12394 29402
rect 12406 29350 12458 29402
rect 12470 29350 12522 29402
rect 23478 29350 23530 29402
rect 23542 29350 23594 29402
rect 23606 29350 23658 29402
rect 23670 29350 23722 29402
rect 23734 29350 23786 29402
rect 1676 29155 1728 29164
rect 1676 29121 1685 29155
rect 1685 29121 1719 29155
rect 1719 29121 1728 29155
rect 1676 29112 1728 29121
rect 33876 29112 33928 29164
rect 34060 29155 34112 29164
rect 34060 29121 34069 29155
rect 34069 29121 34103 29155
rect 34103 29121 34112 29155
rect 34060 29112 34112 29121
rect 1952 28976 2004 29028
rect 34244 29019 34296 29028
rect 34244 28985 34253 29019
rect 34253 28985 34287 29019
rect 34287 28985 34296 29019
rect 34244 28976 34296 28985
rect 34060 28908 34112 28960
rect 6582 28806 6634 28858
rect 6646 28806 6698 28858
rect 6710 28806 6762 28858
rect 6774 28806 6826 28858
rect 6838 28806 6890 28858
rect 17846 28806 17898 28858
rect 17910 28806 17962 28858
rect 17974 28806 18026 28858
rect 18038 28806 18090 28858
rect 18102 28806 18154 28858
rect 29110 28806 29162 28858
rect 29174 28806 29226 28858
rect 29238 28806 29290 28858
rect 29302 28806 29354 28858
rect 29366 28806 29418 28858
rect 33968 28747 34020 28756
rect 33968 28713 33977 28747
rect 33977 28713 34011 28747
rect 34011 28713 34020 28747
rect 33968 28704 34020 28713
rect 12214 28262 12266 28314
rect 12278 28262 12330 28314
rect 12342 28262 12394 28314
rect 12406 28262 12458 28314
rect 12470 28262 12522 28314
rect 23478 28262 23530 28314
rect 23542 28262 23594 28314
rect 23606 28262 23658 28314
rect 23670 28262 23722 28314
rect 23734 28262 23786 28314
rect 20260 28203 20312 28212
rect 20260 28169 20269 28203
rect 20269 28169 20303 28203
rect 20303 28169 20312 28203
rect 20260 28160 20312 28169
rect 1492 27931 1544 27940
rect 1492 27897 1501 27931
rect 1501 27897 1535 27931
rect 1535 27897 1544 27931
rect 1492 27888 1544 27897
rect 30840 28024 30892 28076
rect 34060 28067 34112 28076
rect 34060 28033 34069 28067
rect 34069 28033 34103 28067
rect 34103 28033 34112 28067
rect 34060 28024 34112 28033
rect 34244 27931 34296 27940
rect 34244 27897 34253 27931
rect 34253 27897 34287 27931
rect 34287 27897 34296 27931
rect 34244 27888 34296 27897
rect 2228 27820 2280 27872
rect 34060 27820 34112 27872
rect 6582 27718 6634 27770
rect 6646 27718 6698 27770
rect 6710 27718 6762 27770
rect 6774 27718 6826 27770
rect 6838 27718 6890 27770
rect 17846 27718 17898 27770
rect 17910 27718 17962 27770
rect 17974 27718 18026 27770
rect 18038 27718 18090 27770
rect 18102 27718 18154 27770
rect 29110 27718 29162 27770
rect 29174 27718 29226 27770
rect 29238 27718 29290 27770
rect 29302 27718 29354 27770
rect 29366 27718 29418 27770
rect 19984 27548 20036 27600
rect 6460 27412 6512 27464
rect 20076 27455 20128 27464
rect 20076 27421 20085 27455
rect 20085 27421 20119 27455
rect 20119 27421 20128 27455
rect 20076 27412 20128 27421
rect 20260 27412 20312 27464
rect 20628 27455 20680 27464
rect 20628 27421 20637 27455
rect 20637 27421 20671 27455
rect 20671 27421 20680 27455
rect 20628 27412 20680 27421
rect 18420 27276 18472 27328
rect 21180 27344 21232 27396
rect 20812 27276 20864 27328
rect 21640 27319 21692 27328
rect 21640 27285 21649 27319
rect 21649 27285 21683 27319
rect 21683 27285 21692 27319
rect 21640 27276 21692 27285
rect 12214 27174 12266 27226
rect 12278 27174 12330 27226
rect 12342 27174 12394 27226
rect 12406 27174 12458 27226
rect 12470 27174 12522 27226
rect 23478 27174 23530 27226
rect 23542 27174 23594 27226
rect 23606 27174 23658 27226
rect 23670 27174 23722 27226
rect 23734 27174 23786 27226
rect 18420 27072 18472 27124
rect 18236 26936 18288 26988
rect 19340 27072 19392 27124
rect 20076 27072 20128 27124
rect 19064 26936 19116 26988
rect 19892 26979 19944 26988
rect 16580 26800 16632 26852
rect 19892 26945 19901 26979
rect 19901 26945 19935 26979
rect 19935 26945 19944 26979
rect 19892 26936 19944 26945
rect 19984 26936 20036 26988
rect 20260 26936 20312 26988
rect 21640 27004 21692 27056
rect 21916 26936 21968 26988
rect 20628 26911 20680 26920
rect 20628 26877 20637 26911
rect 20637 26877 20671 26911
rect 20671 26877 20680 26911
rect 20628 26868 20680 26877
rect 24860 27072 24912 27124
rect 34244 26979 34296 26988
rect 34244 26945 34253 26979
rect 34253 26945 34287 26979
rect 34287 26945 34296 26979
rect 34244 26936 34296 26945
rect 20260 26800 20312 26852
rect 18696 26732 18748 26784
rect 20352 26775 20404 26784
rect 20352 26741 20361 26775
rect 20361 26741 20395 26775
rect 20395 26741 20404 26775
rect 20352 26732 20404 26741
rect 21916 26732 21968 26784
rect 32312 26732 32364 26784
rect 34152 26775 34204 26784
rect 34152 26741 34161 26775
rect 34161 26741 34195 26775
rect 34195 26741 34204 26775
rect 34152 26732 34204 26741
rect 6582 26630 6634 26682
rect 6646 26630 6698 26682
rect 6710 26630 6762 26682
rect 6774 26630 6826 26682
rect 6838 26630 6890 26682
rect 17846 26630 17898 26682
rect 17910 26630 17962 26682
rect 17974 26630 18026 26682
rect 18038 26630 18090 26682
rect 18102 26630 18154 26682
rect 29110 26630 29162 26682
rect 29174 26630 29226 26682
rect 29238 26630 29290 26682
rect 29302 26630 29354 26682
rect 29366 26630 29418 26682
rect 18236 26571 18288 26580
rect 18236 26537 18245 26571
rect 18245 26537 18279 26571
rect 18279 26537 18288 26571
rect 18236 26528 18288 26537
rect 21088 26528 21140 26580
rect 21180 26528 21232 26580
rect 3424 26460 3476 26512
rect 2964 26392 3016 26444
rect 1400 26367 1452 26376
rect 1400 26333 1409 26367
rect 1409 26333 1443 26367
rect 1443 26333 1452 26367
rect 1400 26324 1452 26333
rect 18696 26367 18748 26376
rect 18696 26333 18705 26367
rect 18705 26333 18739 26367
rect 18739 26333 18748 26367
rect 18696 26324 18748 26333
rect 19708 26324 19760 26376
rect 20352 26460 20404 26512
rect 32496 26460 32548 26512
rect 21916 26435 21968 26444
rect 20076 26367 20128 26376
rect 20076 26333 20085 26367
rect 20085 26333 20119 26367
rect 20119 26333 20128 26367
rect 20076 26324 20128 26333
rect 20260 26367 20312 26376
rect 20260 26333 20269 26367
rect 20269 26333 20303 26367
rect 20303 26333 20312 26367
rect 21916 26401 21925 26435
rect 21925 26401 21959 26435
rect 21959 26401 21968 26435
rect 21916 26392 21968 26401
rect 20260 26324 20312 26333
rect 20812 26324 20864 26376
rect 21088 26324 21140 26376
rect 31300 26324 31352 26376
rect 34336 26367 34388 26376
rect 34336 26333 34345 26367
rect 34345 26333 34379 26367
rect 34379 26333 34388 26367
rect 34336 26324 34388 26333
rect 20352 26188 20404 26240
rect 20904 26231 20956 26240
rect 20904 26197 20913 26231
rect 20913 26197 20947 26231
rect 20947 26197 20956 26231
rect 20904 26188 20956 26197
rect 21456 26231 21508 26240
rect 21456 26197 21483 26231
rect 21483 26197 21508 26231
rect 21456 26188 21508 26197
rect 12214 26086 12266 26138
rect 12278 26086 12330 26138
rect 12342 26086 12394 26138
rect 12406 26086 12458 26138
rect 12470 26086 12522 26138
rect 23478 26086 23530 26138
rect 23542 26086 23594 26138
rect 23606 26086 23658 26138
rect 23670 26086 23722 26138
rect 23734 26086 23786 26138
rect 19064 25984 19116 26036
rect 19892 25984 19944 26036
rect 17776 25916 17828 25968
rect 18696 25848 18748 25900
rect 19616 25848 19668 25900
rect 19984 25848 20036 25900
rect 20260 25848 20312 25900
rect 20904 25848 20956 25900
rect 21456 25780 21508 25832
rect 25136 25780 25188 25832
rect 20076 25712 20128 25764
rect 18420 25644 18472 25696
rect 20352 25644 20404 25696
rect 20996 25687 21048 25696
rect 20996 25653 21005 25687
rect 21005 25653 21039 25687
rect 21039 25653 21048 25687
rect 20996 25644 21048 25653
rect 6582 25542 6634 25594
rect 6646 25542 6698 25594
rect 6710 25542 6762 25594
rect 6774 25542 6826 25594
rect 6838 25542 6890 25594
rect 17846 25542 17898 25594
rect 17910 25542 17962 25594
rect 17974 25542 18026 25594
rect 18038 25542 18090 25594
rect 18102 25542 18154 25594
rect 29110 25542 29162 25594
rect 29174 25542 29226 25594
rect 29238 25542 29290 25594
rect 29302 25542 29354 25594
rect 29366 25542 29418 25594
rect 19248 25483 19300 25492
rect 19248 25449 19257 25483
rect 19257 25449 19291 25483
rect 19291 25449 19300 25483
rect 19248 25440 19300 25449
rect 19984 25440 20036 25492
rect 20352 25440 20404 25492
rect 18420 25372 18472 25424
rect 33048 25372 33100 25424
rect 19616 25304 19668 25356
rect 20352 25304 20404 25356
rect 9128 25236 9180 25288
rect 19708 25168 19760 25220
rect 6092 25143 6144 25152
rect 6092 25109 6101 25143
rect 6101 25109 6135 25143
rect 6135 25109 6144 25143
rect 6092 25100 6144 25109
rect 20352 25168 20404 25220
rect 20628 25236 20680 25288
rect 20812 25236 20864 25288
rect 34060 25279 34112 25288
rect 34060 25245 34069 25279
rect 34069 25245 34103 25279
rect 34103 25245 34112 25279
rect 34060 25236 34112 25245
rect 31852 25168 31904 25220
rect 20720 25100 20772 25152
rect 20996 25143 21048 25152
rect 20996 25109 21005 25143
rect 21005 25109 21039 25143
rect 21039 25109 21048 25143
rect 20996 25100 21048 25109
rect 34244 25143 34296 25152
rect 34244 25109 34253 25143
rect 34253 25109 34287 25143
rect 34287 25109 34296 25143
rect 34244 25100 34296 25109
rect 12214 24998 12266 25050
rect 12278 24998 12330 25050
rect 12342 24998 12394 25050
rect 12406 24998 12458 25050
rect 12470 24998 12522 25050
rect 23478 24998 23530 25050
rect 23542 24998 23594 25050
rect 23606 24998 23658 25050
rect 23670 24998 23722 25050
rect 23734 24998 23786 25050
rect 20260 24896 20312 24948
rect 2044 24760 2096 24812
rect 34060 24803 34112 24812
rect 34060 24769 34069 24803
rect 34069 24769 34103 24803
rect 34103 24769 34112 24803
rect 34060 24760 34112 24769
rect 1492 24599 1544 24608
rect 1492 24565 1501 24599
rect 1501 24565 1535 24599
rect 1535 24565 1544 24599
rect 1492 24556 1544 24565
rect 2044 24599 2096 24608
rect 2044 24565 2053 24599
rect 2053 24565 2087 24599
rect 2087 24565 2096 24599
rect 2044 24556 2096 24565
rect 20444 24599 20496 24608
rect 20444 24565 20453 24599
rect 20453 24565 20487 24599
rect 20487 24565 20496 24599
rect 20444 24556 20496 24565
rect 34244 24599 34296 24608
rect 34244 24565 34253 24599
rect 34253 24565 34287 24599
rect 34287 24565 34296 24599
rect 34244 24556 34296 24565
rect 6582 24454 6634 24506
rect 6646 24454 6698 24506
rect 6710 24454 6762 24506
rect 6774 24454 6826 24506
rect 6838 24454 6890 24506
rect 17846 24454 17898 24506
rect 17910 24454 17962 24506
rect 17974 24454 18026 24506
rect 18038 24454 18090 24506
rect 18102 24454 18154 24506
rect 29110 24454 29162 24506
rect 29174 24454 29226 24506
rect 29238 24454 29290 24506
rect 29302 24454 29354 24506
rect 29366 24454 29418 24506
rect 16580 24080 16632 24132
rect 33876 24080 33928 24132
rect 34152 24123 34204 24132
rect 34152 24089 34161 24123
rect 34161 24089 34195 24123
rect 34195 24089 34204 24123
rect 34152 24080 34204 24089
rect 1492 24055 1544 24064
rect 1492 24021 1501 24055
rect 1501 24021 1535 24055
rect 1535 24021 1544 24055
rect 1492 24012 1544 24021
rect 20444 24012 20496 24064
rect 12214 23910 12266 23962
rect 12278 23910 12330 23962
rect 12342 23910 12394 23962
rect 12406 23910 12458 23962
rect 12470 23910 12522 23962
rect 23478 23910 23530 23962
rect 23542 23910 23594 23962
rect 23606 23910 23658 23962
rect 23670 23910 23722 23962
rect 23734 23910 23786 23962
rect 34244 23783 34296 23792
rect 34244 23749 34253 23783
rect 34253 23749 34287 23783
rect 34287 23749 34296 23783
rect 34244 23740 34296 23749
rect 4068 23672 4120 23724
rect 20812 23536 20864 23588
rect 1492 23511 1544 23520
rect 1492 23477 1501 23511
rect 1501 23477 1535 23511
rect 1535 23477 1544 23511
rect 1492 23468 1544 23477
rect 6582 23366 6634 23418
rect 6646 23366 6698 23418
rect 6710 23366 6762 23418
rect 6774 23366 6826 23418
rect 6838 23366 6890 23418
rect 17846 23366 17898 23418
rect 17910 23366 17962 23418
rect 17974 23366 18026 23418
rect 18038 23366 18090 23418
rect 18102 23366 18154 23418
rect 29110 23366 29162 23418
rect 29174 23366 29226 23418
rect 29238 23366 29290 23418
rect 29302 23366 29354 23418
rect 29366 23366 29418 23418
rect 33048 23264 33100 23316
rect 34244 23239 34296 23248
rect 34244 23205 34253 23239
rect 34253 23205 34287 23239
rect 34287 23205 34296 23239
rect 34244 23196 34296 23205
rect 12214 22822 12266 22874
rect 12278 22822 12330 22874
rect 12342 22822 12394 22874
rect 12406 22822 12458 22874
rect 12470 22822 12522 22874
rect 23478 22822 23530 22874
rect 23542 22822 23594 22874
rect 23606 22822 23658 22874
rect 23670 22822 23722 22874
rect 23734 22822 23786 22874
rect 6092 22584 6144 22636
rect 31760 22584 31812 22636
rect 31852 22584 31904 22636
rect 34336 22559 34388 22568
rect 34336 22525 34345 22559
rect 34345 22525 34379 22559
rect 34379 22525 34388 22559
rect 34336 22516 34388 22525
rect 1492 22491 1544 22500
rect 1492 22457 1501 22491
rect 1501 22457 1535 22491
rect 1535 22457 1544 22491
rect 1492 22448 1544 22457
rect 2228 22448 2280 22500
rect 6582 22278 6634 22330
rect 6646 22278 6698 22330
rect 6710 22278 6762 22330
rect 6774 22278 6826 22330
rect 6838 22278 6890 22330
rect 17846 22278 17898 22330
rect 17910 22278 17962 22330
rect 17974 22278 18026 22330
rect 18038 22278 18090 22330
rect 18102 22278 18154 22330
rect 29110 22278 29162 22330
rect 29174 22278 29226 22330
rect 29238 22278 29290 22330
rect 29302 22278 29354 22330
rect 29366 22278 29418 22330
rect 34336 22176 34388 22228
rect 34336 21879 34388 21888
rect 34336 21845 34345 21879
rect 34345 21845 34379 21879
rect 34379 21845 34388 21879
rect 34336 21836 34388 21845
rect 12214 21734 12266 21786
rect 12278 21734 12330 21786
rect 12342 21734 12394 21786
rect 12406 21734 12458 21786
rect 12470 21734 12522 21786
rect 23478 21734 23530 21786
rect 23542 21734 23594 21786
rect 23606 21734 23658 21786
rect 23670 21734 23722 21786
rect 23734 21734 23786 21786
rect 1676 21539 1728 21548
rect 1676 21505 1685 21539
rect 1685 21505 1719 21539
rect 1719 21505 1728 21539
rect 1676 21496 1728 21505
rect 31760 21496 31812 21548
rect 34336 21471 34388 21480
rect 34336 21437 34345 21471
rect 34345 21437 34379 21471
rect 34379 21437 34388 21471
rect 34336 21428 34388 21437
rect 1492 21335 1544 21344
rect 1492 21301 1501 21335
rect 1501 21301 1535 21335
rect 1535 21301 1544 21335
rect 1492 21292 1544 21301
rect 6582 21190 6634 21242
rect 6646 21190 6698 21242
rect 6710 21190 6762 21242
rect 6774 21190 6826 21242
rect 6838 21190 6890 21242
rect 17846 21190 17898 21242
rect 17910 21190 17962 21242
rect 17974 21190 18026 21242
rect 18038 21190 18090 21242
rect 18102 21190 18154 21242
rect 29110 21190 29162 21242
rect 29174 21190 29226 21242
rect 29238 21190 29290 21242
rect 29302 21190 29354 21242
rect 29366 21190 29418 21242
rect 33508 20927 33560 20936
rect 33508 20893 33517 20927
rect 33517 20893 33551 20927
rect 33551 20893 33560 20927
rect 33508 20884 33560 20893
rect 2044 20748 2096 20800
rect 12214 20646 12266 20698
rect 12278 20646 12330 20698
rect 12342 20646 12394 20698
rect 12406 20646 12458 20698
rect 12470 20646 12522 20698
rect 23478 20646 23530 20698
rect 23542 20646 23594 20698
rect 23606 20646 23658 20698
rect 23670 20646 23722 20698
rect 23734 20646 23786 20698
rect 34060 20544 34112 20596
rect 34152 20451 34204 20460
rect 34152 20417 34161 20451
rect 34161 20417 34195 20451
rect 34195 20417 34204 20451
rect 34152 20408 34204 20417
rect 1400 20247 1452 20256
rect 1400 20213 1409 20247
rect 1409 20213 1443 20247
rect 1443 20213 1452 20247
rect 1400 20204 1452 20213
rect 6582 20102 6634 20154
rect 6646 20102 6698 20154
rect 6710 20102 6762 20154
rect 6774 20102 6826 20154
rect 6838 20102 6890 20154
rect 17846 20102 17898 20154
rect 17910 20102 17962 20154
rect 17974 20102 18026 20154
rect 18038 20102 18090 20154
rect 18102 20102 18154 20154
rect 29110 20102 29162 20154
rect 29174 20102 29226 20154
rect 29238 20102 29290 20154
rect 29302 20102 29354 20154
rect 29366 20102 29418 20154
rect 34152 20043 34204 20052
rect 34152 20009 34161 20043
rect 34161 20009 34195 20043
rect 34195 20009 34204 20043
rect 34152 20000 34204 20009
rect 1400 19839 1452 19848
rect 1400 19805 1409 19839
rect 1409 19805 1443 19839
rect 1443 19805 1452 19839
rect 1400 19796 1452 19805
rect 34336 19839 34388 19848
rect 34336 19805 34345 19839
rect 34345 19805 34379 19839
rect 34379 19805 34388 19839
rect 34336 19796 34388 19805
rect 17960 19728 18012 19780
rect 12214 19558 12266 19610
rect 12278 19558 12330 19610
rect 12342 19558 12394 19610
rect 12406 19558 12458 19610
rect 12470 19558 12522 19610
rect 23478 19558 23530 19610
rect 23542 19558 23594 19610
rect 23606 19558 23658 19610
rect 23670 19558 23722 19610
rect 23734 19558 23786 19610
rect 1400 19363 1452 19372
rect 1400 19329 1409 19363
rect 1409 19329 1443 19363
rect 1443 19329 1452 19363
rect 1400 19320 1452 19329
rect 31760 19456 31812 19508
rect 17960 19431 18012 19440
rect 17960 19397 17969 19431
rect 17969 19397 18003 19431
rect 18003 19397 18012 19431
rect 17960 19388 18012 19397
rect 20720 19388 20772 19440
rect 18328 19320 18380 19372
rect 34336 19363 34388 19372
rect 34336 19329 34345 19363
rect 34345 19329 34379 19363
rect 34379 19329 34388 19363
rect 34336 19320 34388 19329
rect 28724 19184 28776 19236
rect 17224 19159 17276 19168
rect 17224 19125 17233 19159
rect 17233 19125 17267 19159
rect 17267 19125 17276 19159
rect 17224 19116 17276 19125
rect 19248 19116 19300 19168
rect 6582 19014 6634 19066
rect 6646 19014 6698 19066
rect 6710 19014 6762 19066
rect 6774 19014 6826 19066
rect 6838 19014 6890 19066
rect 17846 19014 17898 19066
rect 17910 19014 17962 19066
rect 17974 19014 18026 19066
rect 18038 19014 18090 19066
rect 18102 19014 18154 19066
rect 29110 19014 29162 19066
rect 29174 19014 29226 19066
rect 29238 19014 29290 19066
rect 29302 19014 29354 19066
rect 29366 19014 29418 19066
rect 2136 18844 2188 18896
rect 12900 18776 12952 18828
rect 2136 18751 2188 18760
rect 2136 18717 2145 18751
rect 2145 18717 2179 18751
rect 2179 18717 2188 18751
rect 2136 18708 2188 18717
rect 2320 18640 2372 18692
rect 17224 18708 17276 18760
rect 29000 18776 29052 18828
rect 33416 18776 33468 18828
rect 18788 18708 18840 18760
rect 20720 18751 20772 18760
rect 20720 18717 20729 18751
rect 20729 18717 20763 18751
rect 20763 18717 20772 18751
rect 20720 18708 20772 18717
rect 29184 18708 29236 18760
rect 34336 18751 34388 18760
rect 34336 18717 34345 18751
rect 34345 18717 34379 18751
rect 34379 18717 34388 18751
rect 34336 18708 34388 18717
rect 1492 18615 1544 18624
rect 1492 18581 1501 18615
rect 1501 18581 1535 18615
rect 1535 18581 1544 18615
rect 1492 18572 1544 18581
rect 1952 18615 2004 18624
rect 1952 18581 1961 18615
rect 1961 18581 1995 18615
rect 1995 18581 2004 18615
rect 1952 18572 2004 18581
rect 2044 18572 2096 18624
rect 18236 18640 18288 18692
rect 18696 18640 18748 18692
rect 22100 18640 22152 18692
rect 31760 18640 31812 18692
rect 19064 18572 19116 18624
rect 19984 18572 20036 18624
rect 20812 18615 20864 18624
rect 20812 18581 20821 18615
rect 20821 18581 20855 18615
rect 20855 18581 20864 18615
rect 20812 18572 20864 18581
rect 29552 18572 29604 18624
rect 12214 18470 12266 18522
rect 12278 18470 12330 18522
rect 12342 18470 12394 18522
rect 12406 18470 12458 18522
rect 12470 18470 12522 18522
rect 23478 18470 23530 18522
rect 23542 18470 23594 18522
rect 23606 18470 23658 18522
rect 23670 18470 23722 18522
rect 23734 18470 23786 18522
rect 1676 18368 1728 18420
rect 3516 18411 3568 18420
rect 3516 18377 3525 18411
rect 3525 18377 3559 18411
rect 3559 18377 3568 18411
rect 3516 18368 3568 18377
rect 4068 18368 4120 18420
rect 12900 18411 12952 18420
rect 12900 18377 12909 18411
rect 12909 18377 12943 18411
rect 12943 18377 12952 18411
rect 12900 18368 12952 18377
rect 16212 18411 16264 18420
rect 16212 18377 16221 18411
rect 16221 18377 16255 18411
rect 16255 18377 16264 18411
rect 16212 18368 16264 18377
rect 1768 18343 1820 18352
rect 1768 18309 1777 18343
rect 1777 18309 1811 18343
rect 1811 18309 1820 18343
rect 1768 18300 1820 18309
rect 3056 18343 3108 18352
rect 3056 18309 3065 18343
rect 3065 18309 3099 18343
rect 3099 18309 3108 18343
rect 3056 18300 3108 18309
rect 3424 18300 3476 18352
rect 6368 18300 6420 18352
rect 6920 18300 6972 18352
rect 8116 18300 8168 18352
rect 29000 18368 29052 18420
rect 29184 18411 29236 18420
rect 29184 18377 29193 18411
rect 29193 18377 29227 18411
rect 29227 18377 29236 18411
rect 29184 18368 29236 18377
rect 29920 18411 29972 18420
rect 29920 18377 29929 18411
rect 29929 18377 29963 18411
rect 29963 18377 29972 18411
rect 29920 18368 29972 18377
rect 30012 18368 30064 18420
rect 31944 18368 31996 18420
rect 19984 18300 20036 18352
rect 24492 18343 24544 18352
rect 24492 18309 24501 18343
rect 24501 18309 24535 18343
rect 24535 18309 24544 18343
rect 24492 18300 24544 18309
rect 27620 18343 27672 18352
rect 27620 18309 27629 18343
rect 27629 18309 27663 18343
rect 27663 18309 27672 18343
rect 27620 18300 27672 18309
rect 29552 18343 29604 18352
rect 29552 18309 29561 18343
rect 29561 18309 29595 18343
rect 29595 18309 29604 18343
rect 29552 18300 29604 18309
rect 31208 18343 31260 18352
rect 31208 18309 31217 18343
rect 31217 18309 31251 18343
rect 31251 18309 31260 18343
rect 31208 18300 31260 18309
rect 32496 18343 32548 18352
rect 32496 18309 32505 18343
rect 32505 18309 32539 18343
rect 32539 18309 32548 18343
rect 32496 18300 32548 18309
rect 1584 18232 1636 18284
rect 3608 18275 3660 18284
rect 3608 18241 3617 18275
rect 3617 18241 3651 18275
rect 3651 18241 3660 18275
rect 3608 18232 3660 18241
rect 6460 18232 6512 18284
rect 7288 18275 7340 18284
rect 7288 18241 7297 18275
rect 7297 18241 7331 18275
rect 7331 18241 7340 18275
rect 7288 18232 7340 18241
rect 15200 18232 15252 18284
rect 15844 18275 15896 18284
rect 15844 18241 15853 18275
rect 15853 18241 15887 18275
rect 15887 18241 15896 18275
rect 15844 18232 15896 18241
rect 16764 18275 16816 18284
rect 16764 18241 16773 18275
rect 16773 18241 16807 18275
rect 16807 18241 16816 18275
rect 16764 18232 16816 18241
rect 17040 18232 17092 18284
rect 19524 18275 19576 18284
rect 1860 18164 1912 18216
rect 19524 18241 19533 18275
rect 19533 18241 19567 18275
rect 19567 18241 19576 18275
rect 19524 18232 19576 18241
rect 19616 18232 19668 18284
rect 2412 18096 2464 18148
rect 1860 18071 1912 18080
rect 1860 18037 1869 18071
rect 1869 18037 1903 18071
rect 1903 18037 1912 18071
rect 1860 18028 1912 18037
rect 2964 18071 3016 18080
rect 2964 18037 2973 18071
rect 2973 18037 3007 18071
rect 3007 18037 3016 18071
rect 2964 18028 3016 18037
rect 6920 18096 6972 18148
rect 16948 18139 17000 18148
rect 16948 18105 16957 18139
rect 16957 18105 16991 18139
rect 16991 18105 17000 18139
rect 16948 18096 17000 18105
rect 17500 18139 17552 18148
rect 17500 18105 17509 18139
rect 17509 18105 17543 18139
rect 17543 18105 17552 18139
rect 17500 18096 17552 18105
rect 16764 18028 16816 18080
rect 19616 18096 19668 18148
rect 18972 18028 19024 18080
rect 22836 18028 22888 18080
rect 25228 18096 25280 18148
rect 27252 18232 27304 18284
rect 29460 18232 29512 18284
rect 30380 18232 30432 18284
rect 32864 18232 32916 18284
rect 33692 18232 33744 18284
rect 34060 18275 34112 18284
rect 34060 18241 34069 18275
rect 34069 18241 34103 18275
rect 34103 18241 34112 18275
rect 34060 18232 34112 18241
rect 30932 18096 30984 18148
rect 30012 18028 30064 18080
rect 30380 18071 30432 18080
rect 30380 18037 30389 18071
rect 30389 18037 30423 18071
rect 30423 18037 30432 18071
rect 30380 18028 30432 18037
rect 31300 18071 31352 18080
rect 31300 18037 31309 18071
rect 31309 18037 31343 18071
rect 31343 18037 31352 18071
rect 31300 18028 31352 18037
rect 33968 18028 34020 18080
rect 34244 18071 34296 18080
rect 34244 18037 34253 18071
rect 34253 18037 34287 18071
rect 34287 18037 34296 18071
rect 34244 18028 34296 18037
rect 6582 17926 6634 17978
rect 6646 17926 6698 17978
rect 6710 17926 6762 17978
rect 6774 17926 6826 17978
rect 6838 17926 6890 17978
rect 17846 17926 17898 17978
rect 17910 17926 17962 17978
rect 17974 17926 18026 17978
rect 18038 17926 18090 17978
rect 18102 17926 18154 17978
rect 29110 17926 29162 17978
rect 29174 17926 29226 17978
rect 29238 17926 29290 17978
rect 29302 17926 29354 17978
rect 29366 17926 29418 17978
rect 2596 17867 2648 17876
rect 2596 17833 2605 17867
rect 2605 17833 2639 17867
rect 2639 17833 2648 17867
rect 2596 17824 2648 17833
rect 15844 17824 15896 17876
rect 16764 17824 16816 17876
rect 16856 17824 16908 17876
rect 17040 17867 17092 17876
rect 17040 17833 17049 17867
rect 17049 17833 17083 17867
rect 17083 17833 17092 17867
rect 17040 17824 17092 17833
rect 18880 17824 18932 17876
rect 32956 17756 33008 17808
rect 1952 17620 2004 17672
rect 17408 17663 17460 17672
rect 17408 17629 17417 17663
rect 17417 17629 17451 17663
rect 17451 17629 17460 17663
rect 17408 17620 17460 17629
rect 2504 17595 2556 17604
rect 2504 17561 2513 17595
rect 2513 17561 2547 17595
rect 2547 17561 2556 17595
rect 2504 17552 2556 17561
rect 8024 17552 8076 17604
rect 32864 17688 32916 17740
rect 27344 17620 27396 17672
rect 17776 17552 17828 17604
rect 18604 17595 18656 17604
rect 18604 17561 18613 17595
rect 18613 17561 18647 17595
rect 18647 17561 18656 17595
rect 18604 17552 18656 17561
rect 19432 17552 19484 17604
rect 32404 17552 32456 17604
rect 2412 17484 2464 17536
rect 17408 17484 17460 17536
rect 25504 17484 25556 17536
rect 12214 17382 12266 17434
rect 12278 17382 12330 17434
rect 12342 17382 12394 17434
rect 12406 17382 12458 17434
rect 12470 17382 12522 17434
rect 23478 17382 23530 17434
rect 23542 17382 23594 17434
rect 23606 17382 23658 17434
rect 23670 17382 23722 17434
rect 23734 17382 23786 17434
rect 17408 17323 17460 17332
rect 17408 17289 17417 17323
rect 17417 17289 17451 17323
rect 17451 17289 17460 17323
rect 17408 17280 17460 17289
rect 25872 17280 25924 17332
rect 19892 17212 19944 17264
rect 34060 17280 34112 17332
rect 17684 17144 17736 17196
rect 29460 17144 29512 17196
rect 29828 17187 29880 17196
rect 29828 17153 29837 17187
rect 29837 17153 29871 17187
rect 29871 17153 29880 17187
rect 29828 17144 29880 17153
rect 33600 17187 33652 17196
rect 33600 17153 33609 17187
rect 33609 17153 33643 17187
rect 33643 17153 33652 17187
rect 33600 17144 33652 17153
rect 18604 17076 18656 17128
rect 33140 17076 33192 17128
rect 1492 17051 1544 17060
rect 1492 17017 1501 17051
rect 1501 17017 1535 17051
rect 1535 17017 1544 17051
rect 1492 17008 1544 17017
rect 34244 17051 34296 17060
rect 34244 17017 34253 17051
rect 34253 17017 34287 17051
rect 34287 17017 34296 17051
rect 34244 17008 34296 17017
rect 6582 16838 6634 16890
rect 6646 16838 6698 16890
rect 6710 16838 6762 16890
rect 6774 16838 6826 16890
rect 6838 16838 6890 16890
rect 17846 16838 17898 16890
rect 17910 16838 17962 16890
rect 17974 16838 18026 16890
rect 18038 16838 18090 16890
rect 18102 16838 18154 16890
rect 29110 16838 29162 16890
rect 29174 16838 29226 16890
rect 29238 16838 29290 16890
rect 29302 16838 29354 16890
rect 29366 16838 29418 16890
rect 17684 16779 17736 16788
rect 17684 16745 17693 16779
rect 17693 16745 17727 16779
rect 17727 16745 17736 16779
rect 17684 16736 17736 16745
rect 34336 16439 34388 16448
rect 34336 16405 34345 16439
rect 34345 16405 34379 16439
rect 34379 16405 34388 16439
rect 34336 16396 34388 16405
rect 12214 16294 12266 16346
rect 12278 16294 12330 16346
rect 12342 16294 12394 16346
rect 12406 16294 12458 16346
rect 12470 16294 12522 16346
rect 23478 16294 23530 16346
rect 23542 16294 23594 16346
rect 23606 16294 23658 16346
rect 23670 16294 23722 16346
rect 23734 16294 23786 16346
rect 18512 16056 18564 16108
rect 31760 15988 31812 16040
rect 34336 16031 34388 16040
rect 34336 15997 34345 16031
rect 34345 15997 34379 16031
rect 34379 15997 34388 16031
rect 34336 15988 34388 15997
rect 1492 15895 1544 15904
rect 1492 15861 1501 15895
rect 1501 15861 1535 15895
rect 1535 15861 1544 15895
rect 1492 15852 1544 15861
rect 6582 15750 6634 15802
rect 6646 15750 6698 15802
rect 6710 15750 6762 15802
rect 6774 15750 6826 15802
rect 6838 15750 6890 15802
rect 17846 15750 17898 15802
rect 17910 15750 17962 15802
rect 17974 15750 18026 15802
rect 18038 15750 18090 15802
rect 18102 15750 18154 15802
rect 29110 15750 29162 15802
rect 29174 15750 29226 15802
rect 29238 15750 29290 15802
rect 29302 15750 29354 15802
rect 29366 15750 29418 15802
rect 2504 15648 2556 15700
rect 1400 15487 1452 15496
rect 1400 15453 1409 15487
rect 1409 15453 1443 15487
rect 1443 15453 1452 15487
rect 1400 15444 1452 15453
rect 34060 15487 34112 15496
rect 34060 15453 34069 15487
rect 34069 15453 34103 15487
rect 34103 15453 34112 15487
rect 34060 15444 34112 15453
rect 34244 15351 34296 15360
rect 34244 15317 34253 15351
rect 34253 15317 34287 15351
rect 34287 15317 34296 15351
rect 34244 15308 34296 15317
rect 12214 15206 12266 15258
rect 12278 15206 12330 15258
rect 12342 15206 12394 15258
rect 12406 15206 12458 15258
rect 12470 15206 12522 15258
rect 23478 15206 23530 15258
rect 23542 15206 23594 15258
rect 23606 15206 23658 15258
rect 23670 15206 23722 15258
rect 23734 15206 23786 15258
rect 18512 15147 18564 15156
rect 18512 15113 18521 15147
rect 18521 15113 18555 15147
rect 18555 15113 18564 15147
rect 18512 15104 18564 15113
rect 34060 15104 34112 15156
rect 31760 15036 31812 15088
rect 18972 14968 19024 15020
rect 34152 15011 34204 15020
rect 34152 14977 34161 15011
rect 34161 14977 34195 15011
rect 34195 14977 34204 15011
rect 34152 14968 34204 14977
rect 11704 14832 11756 14884
rect 18972 14807 19024 14816
rect 18972 14773 18981 14807
rect 18981 14773 19015 14807
rect 19015 14773 19024 14807
rect 18972 14764 19024 14773
rect 6582 14662 6634 14714
rect 6646 14662 6698 14714
rect 6710 14662 6762 14714
rect 6774 14662 6826 14714
rect 6838 14662 6890 14714
rect 17846 14662 17898 14714
rect 17910 14662 17962 14714
rect 17974 14662 18026 14714
rect 18038 14662 18090 14714
rect 18102 14662 18154 14714
rect 29110 14662 29162 14714
rect 29174 14662 29226 14714
rect 29238 14662 29290 14714
rect 29302 14662 29354 14714
rect 29366 14662 29418 14714
rect 34152 14603 34204 14612
rect 34152 14569 34161 14603
rect 34161 14569 34195 14603
rect 34195 14569 34204 14603
rect 34152 14560 34204 14569
rect 11704 14356 11756 14408
rect 34336 14399 34388 14408
rect 34336 14365 34345 14399
rect 34345 14365 34379 14399
rect 34379 14365 34388 14399
rect 34336 14356 34388 14365
rect 1492 14263 1544 14272
rect 1492 14229 1501 14263
rect 1501 14229 1535 14263
rect 1535 14229 1544 14263
rect 1492 14220 1544 14229
rect 34336 14220 34388 14272
rect 12214 14118 12266 14170
rect 12278 14118 12330 14170
rect 12342 14118 12394 14170
rect 12406 14118 12458 14170
rect 12470 14118 12522 14170
rect 23478 14118 23530 14170
rect 23542 14118 23594 14170
rect 23606 14118 23658 14170
rect 23670 14118 23722 14170
rect 23734 14118 23786 14170
rect 33140 13880 33192 13932
rect 34336 13855 34388 13864
rect 34336 13821 34345 13855
rect 34345 13821 34379 13855
rect 34379 13821 34388 13855
rect 34336 13812 34388 13821
rect 6582 13574 6634 13626
rect 6646 13574 6698 13626
rect 6710 13574 6762 13626
rect 6774 13574 6826 13626
rect 6838 13574 6890 13626
rect 17846 13574 17898 13626
rect 17910 13574 17962 13626
rect 17974 13574 18026 13626
rect 18038 13574 18090 13626
rect 18102 13574 18154 13626
rect 29110 13574 29162 13626
rect 29174 13574 29226 13626
rect 29238 13574 29290 13626
rect 29302 13574 29354 13626
rect 29366 13574 29418 13626
rect 1676 13243 1728 13252
rect 1676 13209 1685 13243
rect 1685 13209 1719 13243
rect 1719 13209 1728 13243
rect 1676 13200 1728 13209
rect 17684 13200 17736 13252
rect 33692 13175 33744 13184
rect 33692 13141 33701 13175
rect 33701 13141 33735 13175
rect 33735 13141 33744 13175
rect 33692 13132 33744 13141
rect 34244 13175 34296 13184
rect 34244 13141 34253 13175
rect 34253 13141 34287 13175
rect 34287 13141 34296 13175
rect 34244 13132 34296 13141
rect 12214 13030 12266 13082
rect 12278 13030 12330 13082
rect 12342 13030 12394 13082
rect 12406 13030 12458 13082
rect 12470 13030 12522 13082
rect 23478 13030 23530 13082
rect 23542 13030 23594 13082
rect 23606 13030 23658 13082
rect 23670 13030 23722 13082
rect 23734 13030 23786 13082
rect 2044 12792 2096 12844
rect 17776 12792 17828 12844
rect 1492 12631 1544 12640
rect 1492 12597 1501 12631
rect 1501 12597 1535 12631
rect 1535 12597 1544 12631
rect 1492 12588 1544 12597
rect 2044 12631 2096 12640
rect 2044 12597 2053 12631
rect 2053 12597 2087 12631
rect 2087 12597 2096 12631
rect 2044 12588 2096 12597
rect 34244 12631 34296 12640
rect 34244 12597 34253 12631
rect 34253 12597 34287 12631
rect 34287 12597 34296 12631
rect 34244 12588 34296 12597
rect 6582 12486 6634 12538
rect 6646 12486 6698 12538
rect 6710 12486 6762 12538
rect 6774 12486 6826 12538
rect 6838 12486 6890 12538
rect 17846 12486 17898 12538
rect 17910 12486 17962 12538
rect 17974 12486 18026 12538
rect 18038 12486 18090 12538
rect 18102 12486 18154 12538
rect 29110 12486 29162 12538
rect 29174 12486 29226 12538
rect 29238 12486 29290 12538
rect 29302 12486 29354 12538
rect 29366 12486 29418 12538
rect 12214 11942 12266 11994
rect 12278 11942 12330 11994
rect 12342 11942 12394 11994
rect 12406 11942 12458 11994
rect 12470 11942 12522 11994
rect 23478 11942 23530 11994
rect 23542 11942 23594 11994
rect 23606 11942 23658 11994
rect 23670 11942 23722 11994
rect 23734 11942 23786 11994
rect 1400 11679 1452 11688
rect 1400 11645 1409 11679
rect 1409 11645 1443 11679
rect 1443 11645 1452 11679
rect 1400 11636 1452 11645
rect 18880 11568 18932 11620
rect 19248 11568 19300 11620
rect 34244 11611 34296 11620
rect 34244 11577 34253 11611
rect 34253 11577 34287 11611
rect 34287 11577 34296 11611
rect 34244 11568 34296 11577
rect 6582 11398 6634 11450
rect 6646 11398 6698 11450
rect 6710 11398 6762 11450
rect 6774 11398 6826 11450
rect 6838 11398 6890 11450
rect 17846 11398 17898 11450
rect 17910 11398 17962 11450
rect 17974 11398 18026 11450
rect 18038 11398 18090 11450
rect 18102 11398 18154 11450
rect 29110 11398 29162 11450
rect 29174 11398 29226 11450
rect 29238 11398 29290 11450
rect 29302 11398 29354 11450
rect 29366 11398 29418 11450
rect 1400 11339 1452 11348
rect 1400 11305 1409 11339
rect 1409 11305 1443 11339
rect 1443 11305 1452 11339
rect 1400 11296 1452 11305
rect 12214 10854 12266 10906
rect 12278 10854 12330 10906
rect 12342 10854 12394 10906
rect 12406 10854 12458 10906
rect 12470 10854 12522 10906
rect 23478 10854 23530 10906
rect 23542 10854 23594 10906
rect 23606 10854 23658 10906
rect 23670 10854 23722 10906
rect 23734 10854 23786 10906
rect 1584 10795 1636 10804
rect 1584 10761 1593 10795
rect 1593 10761 1627 10795
rect 1627 10761 1636 10795
rect 1584 10752 1636 10761
rect 1400 10659 1452 10668
rect 1400 10625 1409 10659
rect 1409 10625 1443 10659
rect 1443 10625 1452 10659
rect 1400 10616 1452 10625
rect 6582 10310 6634 10362
rect 6646 10310 6698 10362
rect 6710 10310 6762 10362
rect 6774 10310 6826 10362
rect 6838 10310 6890 10362
rect 17846 10310 17898 10362
rect 17910 10310 17962 10362
rect 17974 10310 18026 10362
rect 18038 10310 18090 10362
rect 18102 10310 18154 10362
rect 29110 10310 29162 10362
rect 29174 10310 29226 10362
rect 29238 10310 29290 10362
rect 29302 10310 29354 10362
rect 29366 10310 29418 10362
rect 33600 10208 33652 10260
rect 34336 10047 34388 10056
rect 34336 10013 34345 10047
rect 34345 10013 34379 10047
rect 34379 10013 34388 10047
rect 34336 10004 34388 10013
rect 17316 9936 17368 9988
rect 33692 9868 33744 9920
rect 12214 9766 12266 9818
rect 12278 9766 12330 9818
rect 12342 9766 12394 9818
rect 12406 9766 12458 9818
rect 12470 9766 12522 9818
rect 23478 9766 23530 9818
rect 23542 9766 23594 9818
rect 23606 9766 23658 9818
rect 23670 9766 23722 9818
rect 23734 9766 23786 9818
rect 18512 9528 18564 9580
rect 2044 9324 2096 9376
rect 18512 9367 18564 9376
rect 18512 9333 18521 9367
rect 18521 9333 18555 9367
rect 18555 9333 18564 9367
rect 18512 9324 18564 9333
rect 6582 9222 6634 9274
rect 6646 9222 6698 9274
rect 6710 9222 6762 9274
rect 6774 9222 6826 9274
rect 6838 9222 6890 9274
rect 17846 9222 17898 9274
rect 17910 9222 17962 9274
rect 17974 9222 18026 9274
rect 18038 9222 18090 9274
rect 18102 9222 18154 9274
rect 29110 9222 29162 9274
rect 29174 9222 29226 9274
rect 29238 9222 29290 9274
rect 29302 9222 29354 9274
rect 29366 9222 29418 9274
rect 18236 8916 18288 8968
rect 19340 8848 19392 8900
rect 1492 8823 1544 8832
rect 1492 8789 1501 8823
rect 1501 8789 1535 8823
rect 1535 8789 1544 8823
rect 1492 8780 1544 8789
rect 34244 8823 34296 8832
rect 34244 8789 34253 8823
rect 34253 8789 34287 8823
rect 34287 8789 34296 8823
rect 34244 8780 34296 8789
rect 12214 8678 12266 8730
rect 12278 8678 12330 8730
rect 12342 8678 12394 8730
rect 12406 8678 12458 8730
rect 12470 8678 12522 8730
rect 23478 8678 23530 8730
rect 23542 8678 23594 8730
rect 23606 8678 23658 8730
rect 23670 8678 23722 8730
rect 23734 8678 23786 8730
rect 34244 8483 34296 8492
rect 34244 8449 34253 8483
rect 34253 8449 34287 8483
rect 34287 8449 34296 8483
rect 34244 8440 34296 8449
rect 18972 8304 19024 8356
rect 6582 8134 6634 8186
rect 6646 8134 6698 8186
rect 6710 8134 6762 8186
rect 6774 8134 6826 8186
rect 6838 8134 6890 8186
rect 17846 8134 17898 8186
rect 17910 8134 17962 8186
rect 17974 8134 18026 8186
rect 18038 8134 18090 8186
rect 18102 8134 18154 8186
rect 29110 8134 29162 8186
rect 29174 8134 29226 8186
rect 29238 8134 29290 8186
rect 29302 8134 29354 8186
rect 29366 8134 29418 8186
rect 10968 7828 11020 7880
rect 33968 7828 34020 7880
rect 1492 7735 1544 7744
rect 1492 7701 1501 7735
rect 1501 7701 1535 7735
rect 1535 7701 1544 7735
rect 1492 7692 1544 7701
rect 34244 7735 34296 7744
rect 34244 7701 34253 7735
rect 34253 7701 34287 7735
rect 34287 7701 34296 7735
rect 34244 7692 34296 7701
rect 12214 7590 12266 7642
rect 12278 7590 12330 7642
rect 12342 7590 12394 7642
rect 12406 7590 12458 7642
rect 12470 7590 12522 7642
rect 23478 7590 23530 7642
rect 23542 7590 23594 7642
rect 23606 7590 23658 7642
rect 23670 7590 23722 7642
rect 23734 7590 23786 7642
rect 2044 7352 2096 7404
rect 32404 7352 32456 7404
rect 1492 7191 1544 7200
rect 1492 7157 1501 7191
rect 1501 7157 1535 7191
rect 1535 7157 1544 7191
rect 1492 7148 1544 7157
rect 2044 7191 2096 7200
rect 2044 7157 2053 7191
rect 2053 7157 2087 7191
rect 2087 7157 2096 7191
rect 2044 7148 2096 7157
rect 34244 7191 34296 7200
rect 34244 7157 34253 7191
rect 34253 7157 34287 7191
rect 34287 7157 34296 7191
rect 34244 7148 34296 7157
rect 6582 7046 6634 7098
rect 6646 7046 6698 7098
rect 6710 7046 6762 7098
rect 6774 7046 6826 7098
rect 6838 7046 6890 7098
rect 17846 7046 17898 7098
rect 17910 7046 17962 7098
rect 17974 7046 18026 7098
rect 18038 7046 18090 7098
rect 18102 7046 18154 7098
rect 29110 7046 29162 7098
rect 29174 7046 29226 7098
rect 29238 7046 29290 7098
rect 29302 7046 29354 7098
rect 29366 7046 29418 7098
rect 12214 6502 12266 6554
rect 12278 6502 12330 6554
rect 12342 6502 12394 6554
rect 12406 6502 12458 6554
rect 12470 6502 12522 6554
rect 23478 6502 23530 6554
rect 23542 6502 23594 6554
rect 23606 6502 23658 6554
rect 23670 6502 23722 6554
rect 23734 6502 23786 6554
rect 2964 6264 3016 6316
rect 34244 6307 34296 6316
rect 34244 6273 34253 6307
rect 34253 6273 34287 6307
rect 34287 6273 34296 6307
rect 34244 6264 34296 6273
rect 1492 6171 1544 6180
rect 1492 6137 1501 6171
rect 1501 6137 1535 6171
rect 1535 6137 1544 6171
rect 1492 6128 1544 6137
rect 19984 6060 20036 6112
rect 6582 5958 6634 6010
rect 6646 5958 6698 6010
rect 6710 5958 6762 6010
rect 6774 5958 6826 6010
rect 6838 5958 6890 6010
rect 17846 5958 17898 6010
rect 17910 5958 17962 6010
rect 17974 5958 18026 6010
rect 18038 5958 18090 6010
rect 18102 5958 18154 6010
rect 29110 5958 29162 6010
rect 29174 5958 29226 6010
rect 29238 5958 29290 6010
rect 29302 5958 29354 6010
rect 29366 5958 29418 6010
rect 34336 5559 34388 5568
rect 34336 5525 34345 5559
rect 34345 5525 34379 5559
rect 34379 5525 34388 5559
rect 34336 5516 34388 5525
rect 12214 5414 12266 5466
rect 12278 5414 12330 5466
rect 12342 5414 12394 5466
rect 12406 5414 12458 5466
rect 12470 5414 12522 5466
rect 23478 5414 23530 5466
rect 23542 5414 23594 5466
rect 23606 5414 23658 5466
rect 23670 5414 23722 5466
rect 23734 5414 23786 5466
rect 10968 5355 11020 5364
rect 10968 5321 10977 5355
rect 10977 5321 11011 5355
rect 11011 5321 11020 5355
rect 10968 5312 11020 5321
rect 13636 5176 13688 5228
rect 17776 5108 17828 5160
rect 30104 5108 30156 5160
rect 34336 5151 34388 5160
rect 34336 5117 34345 5151
rect 34345 5117 34379 5151
rect 34379 5117 34388 5151
rect 34336 5108 34388 5117
rect 1492 5015 1544 5024
rect 1492 4981 1501 5015
rect 1501 4981 1535 5015
rect 1535 4981 1544 5015
rect 1492 4972 1544 4981
rect 6582 4870 6634 4922
rect 6646 4870 6698 4922
rect 6710 4870 6762 4922
rect 6774 4870 6826 4922
rect 6838 4870 6890 4922
rect 17846 4870 17898 4922
rect 17910 4870 17962 4922
rect 17974 4870 18026 4922
rect 18038 4870 18090 4922
rect 18102 4870 18154 4922
rect 29110 4870 29162 4922
rect 29174 4870 29226 4922
rect 29238 4870 29290 4922
rect 29302 4870 29354 4922
rect 29366 4870 29418 4922
rect 17776 4700 17828 4752
rect 1400 4471 1452 4480
rect 1400 4437 1409 4471
rect 1409 4437 1443 4471
rect 1443 4437 1452 4471
rect 1400 4428 1452 4437
rect 2044 4428 2096 4480
rect 30104 4632 30156 4684
rect 20352 4496 20404 4548
rect 17592 4428 17644 4480
rect 34244 4471 34296 4480
rect 34244 4437 34253 4471
rect 34253 4437 34287 4471
rect 34287 4437 34296 4471
rect 34244 4428 34296 4437
rect 12214 4326 12266 4378
rect 12278 4326 12330 4378
rect 12342 4326 12394 4378
rect 12406 4326 12458 4378
rect 12470 4326 12522 4378
rect 23478 4326 23530 4378
rect 23542 4326 23594 4378
rect 23606 4326 23658 4378
rect 23670 4326 23722 4378
rect 23734 4326 23786 4378
rect 1400 4131 1452 4140
rect 1400 4097 1409 4131
rect 1409 4097 1443 4131
rect 1443 4097 1452 4131
rect 1400 4088 1452 4097
rect 3056 4088 3108 4140
rect 33876 4088 33928 4140
rect 11612 3952 11664 4004
rect 2044 3927 2096 3936
rect 2044 3893 2053 3927
rect 2053 3893 2087 3927
rect 2087 3893 2096 3927
rect 2044 3884 2096 3893
rect 3056 3884 3108 3936
rect 33876 3884 33928 3936
rect 34244 3927 34296 3936
rect 34244 3893 34253 3927
rect 34253 3893 34287 3927
rect 34287 3893 34296 3927
rect 34244 3884 34296 3893
rect 6582 3782 6634 3834
rect 6646 3782 6698 3834
rect 6710 3782 6762 3834
rect 6774 3782 6826 3834
rect 6838 3782 6890 3834
rect 17846 3782 17898 3834
rect 17910 3782 17962 3834
rect 17974 3782 18026 3834
rect 18038 3782 18090 3834
rect 18102 3782 18154 3834
rect 29110 3782 29162 3834
rect 29174 3782 29226 3834
rect 29238 3782 29290 3834
rect 29302 3782 29354 3834
rect 29366 3782 29418 3834
rect 8116 3723 8168 3732
rect 8116 3689 8125 3723
rect 8125 3689 8159 3723
rect 8159 3689 8168 3723
rect 8116 3680 8168 3689
rect 14556 3680 14608 3732
rect 20 3612 72 3664
rect 6828 3612 6880 3664
rect 13728 3612 13780 3664
rect 4436 3544 4488 3596
rect 17408 3612 17460 3664
rect 20536 3680 20588 3732
rect 34520 3680 34572 3732
rect 18512 3612 18564 3664
rect 17132 3544 17184 3596
rect 34796 3612 34848 3664
rect 1860 3476 1912 3528
rect 2044 3476 2096 3528
rect 16672 3519 16724 3528
rect 16672 3485 16681 3519
rect 16681 3485 16715 3519
rect 16715 3485 16724 3519
rect 16672 3476 16724 3485
rect 17224 3476 17276 3528
rect 29736 3476 29788 3528
rect 31852 3476 31904 3528
rect 32404 3519 32456 3528
rect 32404 3485 32413 3519
rect 32413 3485 32447 3519
rect 32447 3485 32456 3519
rect 32404 3476 32456 3485
rect 4252 3408 4304 3460
rect 17776 3408 17828 3460
rect 19156 3408 19208 3460
rect 19708 3408 19760 3460
rect 34520 3408 34572 3460
rect 35440 3408 35492 3460
rect 664 3340 716 3392
rect 2964 3383 3016 3392
rect 2964 3349 2973 3383
rect 2973 3349 3007 3383
rect 3007 3349 3016 3383
rect 2964 3340 3016 3349
rect 3792 3383 3844 3392
rect 3792 3349 3801 3383
rect 3801 3349 3835 3383
rect 3835 3349 3844 3383
rect 3792 3340 3844 3349
rect 4160 3383 4212 3392
rect 4160 3349 4169 3383
rect 4169 3349 4203 3383
rect 4203 3349 4212 3383
rect 4160 3340 4212 3349
rect 11704 3340 11756 3392
rect 17500 3340 17552 3392
rect 18880 3340 18932 3392
rect 33140 3383 33192 3392
rect 33140 3349 33149 3383
rect 33149 3349 33183 3383
rect 33183 3349 33192 3383
rect 33140 3340 33192 3349
rect 12214 3238 12266 3290
rect 12278 3238 12330 3290
rect 12342 3238 12394 3290
rect 12406 3238 12458 3290
rect 12470 3238 12522 3290
rect 23478 3238 23530 3290
rect 23542 3238 23594 3290
rect 23606 3238 23658 3290
rect 23670 3238 23722 3290
rect 23734 3238 23786 3290
rect 13636 3179 13688 3188
rect 4436 3068 4488 3120
rect 2412 3000 2464 3052
rect 4252 3043 4304 3052
rect 4252 3009 4261 3043
rect 4261 3009 4295 3043
rect 4295 3009 4304 3043
rect 4252 3000 4304 3009
rect 6828 3043 6880 3052
rect 6828 3009 6837 3043
rect 6837 3009 6871 3043
rect 6871 3009 6880 3043
rect 6828 3000 6880 3009
rect 7748 3000 7800 3052
rect 13636 3145 13645 3179
rect 13645 3145 13679 3179
rect 13679 3145 13688 3179
rect 13636 3136 13688 3145
rect 13728 3136 13780 3188
rect 17776 3068 17828 3120
rect 19708 3136 19760 3188
rect 20352 3136 20404 3188
rect 22836 3179 22888 3188
rect 22836 3145 22845 3179
rect 22845 3145 22879 3179
rect 22879 3145 22888 3179
rect 22836 3136 22888 3145
rect 25136 3179 25188 3188
rect 25136 3145 25145 3179
rect 25145 3145 25179 3179
rect 25179 3145 25188 3179
rect 25136 3136 25188 3145
rect 29736 3179 29788 3188
rect 29736 3145 29745 3179
rect 29745 3145 29779 3179
rect 29779 3145 29788 3179
rect 29736 3136 29788 3145
rect 11612 3043 11664 3052
rect 2964 2932 3016 2984
rect 11612 3009 11621 3043
rect 11621 3009 11655 3043
rect 11655 3009 11664 3043
rect 11612 3000 11664 3009
rect 13544 3000 13596 3052
rect 14372 3043 14424 3052
rect 14372 3009 14381 3043
rect 14381 3009 14415 3043
rect 14415 3009 14424 3043
rect 14372 3000 14424 3009
rect 17132 3043 17184 3052
rect 17132 3009 17141 3043
rect 17141 3009 17175 3043
rect 17175 3009 17184 3043
rect 17132 3000 17184 3009
rect 17408 3043 17460 3052
rect 17408 3009 17417 3043
rect 17417 3009 17451 3043
rect 17451 3009 17460 3043
rect 17408 3000 17460 3009
rect 18328 3000 18380 3052
rect 18512 3043 18564 3052
rect 18512 3009 18521 3043
rect 18521 3009 18555 3043
rect 18555 3009 18564 3043
rect 18512 3000 18564 3009
rect 28632 3068 28684 3120
rect 30380 3068 30432 3120
rect 11704 2932 11756 2984
rect 19248 2932 19300 2984
rect 2596 2864 2648 2916
rect 10232 2864 10284 2916
rect 10968 2864 11020 2916
rect 12440 2864 12492 2916
rect 21824 3000 21876 3052
rect 21916 3000 21968 3052
rect 25136 3000 25188 3052
rect 25504 3000 25556 3052
rect 29644 3000 29696 3052
rect 31300 3000 31352 3052
rect 32404 3000 32456 3052
rect 1952 2796 2004 2848
rect 2872 2796 2924 2848
rect 3884 2796 3936 2848
rect 4528 2796 4580 2848
rect 5816 2796 5868 2848
rect 6460 2796 6512 2848
rect 9036 2796 9088 2848
rect 12992 2796 13044 2848
rect 13544 2796 13596 2848
rect 13728 2796 13780 2848
rect 15200 2796 15252 2848
rect 19340 2796 19392 2848
rect 28080 2932 28132 2984
rect 33508 2975 33560 2984
rect 33508 2941 33517 2975
rect 33517 2941 33551 2975
rect 33551 2941 33560 2975
rect 33508 2932 33560 2941
rect 20812 2864 20864 2916
rect 32404 2864 32456 2916
rect 24492 2796 24544 2848
rect 27068 2796 27120 2848
rect 29460 2839 29512 2848
rect 29460 2805 29469 2839
rect 29469 2805 29503 2839
rect 29503 2805 29512 2839
rect 29460 2796 29512 2805
rect 32220 2796 32272 2848
rect 32864 2796 32916 2848
rect 6582 2694 6634 2746
rect 6646 2694 6698 2746
rect 6710 2694 6762 2746
rect 6774 2694 6826 2746
rect 6838 2694 6890 2746
rect 17846 2694 17898 2746
rect 17910 2694 17962 2746
rect 17974 2694 18026 2746
rect 18038 2694 18090 2746
rect 18102 2694 18154 2746
rect 29110 2694 29162 2746
rect 29174 2694 29226 2746
rect 29238 2694 29290 2746
rect 29302 2694 29354 2746
rect 29366 2694 29418 2746
rect 14372 2592 14424 2644
rect 17316 2592 17368 2644
rect 18328 2592 18380 2644
rect 1400 2456 1452 2508
rect 2596 2456 2648 2508
rect 2504 2388 2556 2440
rect 3240 2388 3292 2440
rect 4160 2524 4212 2576
rect 6368 2524 6420 2576
rect 3608 2456 3660 2508
rect 7288 2456 7340 2508
rect 3424 2388 3476 2440
rect 3792 2431 3844 2440
rect 3792 2397 3801 2431
rect 3801 2397 3835 2431
rect 3835 2397 3844 2431
rect 3792 2388 3844 2397
rect 2872 2320 2924 2372
rect 4528 2388 4580 2440
rect 5816 2388 5868 2440
rect 8024 2388 8076 2440
rect 8116 2388 8168 2440
rect 9036 2388 9088 2440
rect 10232 2431 10284 2440
rect 10232 2397 10241 2431
rect 10241 2397 10275 2431
rect 10275 2397 10284 2431
rect 10232 2388 10284 2397
rect 10968 2431 11020 2440
rect 10968 2397 10977 2431
rect 10977 2397 11011 2431
rect 11011 2397 11020 2431
rect 10968 2388 11020 2397
rect 12440 2388 12492 2440
rect 14556 2524 14608 2576
rect 12992 2456 13044 2508
rect 19432 2524 19484 2576
rect 21824 2592 21876 2644
rect 28632 2635 28684 2644
rect 28632 2601 28641 2635
rect 28641 2601 28675 2635
rect 28675 2601 28684 2635
rect 28632 2592 28684 2601
rect 32956 2567 33008 2576
rect 32956 2533 32965 2567
rect 32965 2533 32999 2567
rect 32999 2533 33008 2567
rect 32956 2524 33008 2533
rect 13728 2431 13780 2440
rect 11888 2320 11940 2372
rect 13728 2397 13737 2431
rect 13737 2397 13771 2431
rect 13771 2397 13780 2431
rect 13728 2388 13780 2397
rect 18696 2456 18748 2508
rect 19156 2456 19208 2508
rect 19524 2499 19576 2508
rect 19524 2465 19533 2499
rect 19533 2465 19567 2499
rect 19567 2465 19576 2499
rect 19524 2456 19576 2465
rect 20536 2456 20588 2508
rect 27252 2499 27304 2508
rect 14832 2388 14884 2440
rect 16764 2388 16816 2440
rect 16948 2431 17000 2440
rect 16948 2397 16957 2431
rect 16957 2397 16991 2431
rect 16991 2397 17000 2431
rect 16948 2388 17000 2397
rect 17500 2431 17552 2440
rect 17500 2397 17509 2431
rect 17509 2397 17543 2431
rect 17543 2397 17552 2431
rect 17500 2388 17552 2397
rect 18052 2388 18104 2440
rect 18880 2431 18932 2440
rect 18880 2397 18889 2431
rect 18889 2397 18923 2431
rect 18923 2397 18932 2431
rect 18880 2388 18932 2397
rect 22100 2431 22152 2440
rect 16856 2320 16908 2372
rect 18788 2320 18840 2372
rect 22100 2397 22109 2431
rect 22109 2397 22143 2431
rect 22143 2397 22152 2431
rect 22100 2388 22152 2397
rect 22836 2388 22888 2440
rect 23480 2431 23532 2440
rect 23480 2397 23489 2431
rect 23489 2397 23523 2431
rect 23523 2397 23532 2431
rect 27252 2465 27261 2499
rect 27261 2465 27295 2499
rect 27295 2465 27304 2499
rect 27252 2456 27304 2465
rect 29828 2499 29880 2508
rect 29828 2465 29837 2499
rect 29837 2465 29871 2499
rect 29871 2465 29880 2499
rect 29828 2456 29880 2465
rect 31852 2456 31904 2508
rect 23480 2388 23532 2397
rect 25228 2431 25280 2440
rect 25228 2397 25237 2431
rect 25237 2397 25271 2431
rect 25271 2397 25280 2431
rect 25228 2388 25280 2397
rect 2780 2252 2832 2304
rect 7104 2252 7156 2304
rect 8392 2252 8444 2304
rect 9680 2252 9732 2304
rect 11152 2295 11204 2304
rect 11152 2261 11161 2295
rect 11161 2261 11195 2295
rect 11195 2261 11204 2295
rect 11152 2252 11204 2261
rect 11612 2252 11664 2304
rect 12072 2252 12124 2304
rect 12900 2252 12952 2304
rect 13728 2252 13780 2304
rect 14188 2252 14240 2304
rect 16120 2252 16172 2304
rect 17408 2252 17460 2304
rect 19984 2252 20036 2304
rect 21272 2252 21324 2304
rect 22560 2252 22612 2304
rect 23848 2252 23900 2304
rect 25136 2252 25188 2304
rect 26424 2252 26476 2304
rect 28080 2431 28132 2440
rect 28080 2397 28089 2431
rect 28089 2397 28123 2431
rect 28123 2397 28132 2431
rect 28080 2388 28132 2397
rect 28356 2388 28408 2440
rect 29000 2388 29052 2440
rect 29460 2388 29512 2440
rect 30932 2431 30984 2440
rect 30932 2397 30941 2431
rect 30941 2397 30975 2431
rect 30975 2397 30984 2431
rect 30932 2388 30984 2397
rect 31576 2388 31628 2440
rect 32404 2431 32456 2440
rect 32404 2397 32413 2431
rect 32413 2397 32447 2431
rect 32447 2397 32456 2431
rect 32404 2388 32456 2397
rect 33876 2456 33928 2508
rect 33140 2363 33192 2372
rect 33140 2329 33149 2363
rect 33149 2329 33183 2363
rect 33183 2329 33192 2363
rect 33140 2320 33192 2329
rect 27712 2252 27764 2304
rect 30288 2252 30340 2304
rect 32588 2295 32640 2304
rect 32588 2261 32597 2295
rect 32597 2261 32631 2295
rect 32631 2261 32640 2295
rect 32588 2252 32640 2261
rect 12214 2150 12266 2202
rect 12278 2150 12330 2202
rect 12342 2150 12394 2202
rect 12406 2150 12458 2202
rect 12470 2150 12522 2202
rect 23478 2150 23530 2202
rect 23542 2150 23594 2202
rect 23606 2150 23658 2202
rect 23670 2150 23722 2202
rect 23734 2150 23786 2202
rect 2504 2048 2556 2100
rect 3240 1980 3292 2032
rect 11888 2048 11940 2100
rect 17224 2048 17276 2100
rect 16672 1980 16724 2032
rect 11152 1912 11204 1964
rect 18512 1912 18564 1964
rect 18236 1844 18288 1896
rect 8024 1776 8076 1828
rect 15200 1776 15252 1828
<< metal2 >>
rect 18 35200 74 36000
rect 662 35306 718 36000
rect 662 35278 1072 35306
rect 662 35200 718 35278
rect 32 32910 60 35200
rect 1044 33522 1072 35278
rect 1306 35200 1362 36000
rect 2594 35306 2650 36000
rect 2962 35456 3018 35465
rect 2962 35391 3018 35400
rect 2594 35278 2728 35306
rect 2594 35200 2650 35278
rect 1032 33516 1084 33522
rect 1032 33458 1084 33464
rect 1320 33046 1348 35200
rect 2134 34096 2190 34105
rect 2700 34082 2728 35278
rect 2870 34776 2926 34785
rect 2870 34711 2926 34720
rect 2700 34054 2820 34082
rect 2134 34031 2190 34040
rect 1308 33040 1360 33046
rect 1308 32982 1360 32988
rect 2148 32910 2176 34031
rect 2792 33590 2820 34054
rect 2780 33584 2832 33590
rect 2780 33526 2832 33532
rect 2228 33516 2280 33522
rect 2228 33458 2280 33464
rect 2240 33114 2268 33458
rect 2596 33312 2648 33318
rect 2596 33254 2648 33260
rect 2228 33108 2280 33114
rect 2228 33050 2280 33056
rect 20 32904 72 32910
rect 20 32846 72 32852
rect 1308 32904 1360 32910
rect 1308 32846 1360 32852
rect 2136 32904 2188 32910
rect 2136 32846 2188 32852
rect 1320 32502 1348 32846
rect 1860 32836 1912 32842
rect 1860 32778 1912 32784
rect 1308 32496 1360 32502
rect 1308 32438 1360 32444
rect 1400 32360 1452 32366
rect 1400 32302 1452 32308
rect 1768 32360 1820 32366
rect 1768 32302 1820 32308
rect 1412 32065 1440 32302
rect 1398 32056 1454 32065
rect 1398 31991 1454 32000
rect 1412 31482 1440 31991
rect 1674 31920 1730 31929
rect 1674 31855 1730 31864
rect 1688 31822 1716 31855
rect 1676 31816 1728 31822
rect 1676 31758 1728 31764
rect 1492 31680 1544 31686
rect 1492 31622 1544 31628
rect 1400 31476 1452 31482
rect 1400 31418 1452 31424
rect 1504 31385 1532 31622
rect 1490 31376 1546 31385
rect 1490 31311 1546 31320
rect 1490 30696 1546 30705
rect 1490 30631 1546 30640
rect 1504 30598 1532 30631
rect 1492 30592 1544 30598
rect 1492 30534 1544 30540
rect 1492 29504 1544 29510
rect 1492 29446 1544 29452
rect 1504 29345 1532 29446
rect 1490 29336 1546 29345
rect 1490 29271 1546 29280
rect 1676 29164 1728 29170
rect 1676 29106 1728 29112
rect 1688 28665 1716 29106
rect 1674 28656 1730 28665
rect 1674 28591 1730 28600
rect 1490 27976 1546 27985
rect 1490 27911 1492 27920
rect 1544 27911 1546 27920
rect 1492 27882 1544 27888
rect 1400 26376 1452 26382
rect 1400 26318 1452 26324
rect 1412 25945 1440 26318
rect 1398 25936 1454 25945
rect 1398 25871 1454 25880
rect 1492 24608 1544 24614
rect 1490 24576 1492 24585
rect 1544 24576 1546 24585
rect 1490 24511 1546 24520
rect 1492 24064 1544 24070
rect 1492 24006 1544 24012
rect 1504 23905 1532 24006
rect 1490 23896 1546 23905
rect 1490 23831 1546 23840
rect 1492 23520 1544 23526
rect 1492 23462 1544 23468
rect 1504 23225 1532 23462
rect 1490 23216 1546 23225
rect 1490 23151 1546 23160
rect 1490 22536 1546 22545
rect 1490 22471 1492 22480
rect 1544 22471 1546 22480
rect 1492 22442 1544 22448
rect 1676 21548 1728 21554
rect 1676 21490 1728 21496
rect 1492 21344 1544 21350
rect 1492 21286 1544 21292
rect 1504 21185 1532 21286
rect 1490 21176 1546 21185
rect 1490 21111 1546 21120
rect 1400 20256 1452 20262
rect 1400 20198 1452 20204
rect 1412 19854 1440 20198
rect 1400 19848 1452 19854
rect 1398 19816 1400 19825
rect 1452 19816 1454 19825
rect 1398 19751 1454 19760
rect 1400 19372 1452 19378
rect 1400 19314 1452 19320
rect 1412 19145 1440 19314
rect 1398 19136 1454 19145
rect 1398 19071 1454 19080
rect 1492 18624 1544 18630
rect 1492 18566 1544 18572
rect 1504 17785 1532 18566
rect 1688 18426 1716 21490
rect 1676 18420 1728 18426
rect 1676 18362 1728 18368
rect 1780 18358 1808 32302
rect 1768 18352 1820 18358
rect 1768 18294 1820 18300
rect 1584 18284 1636 18290
rect 1584 18226 1636 18232
rect 1490 17776 1546 17785
rect 1490 17711 1546 17720
rect 1490 17096 1546 17105
rect 1490 17031 1492 17040
rect 1544 17031 1546 17040
rect 1492 17002 1544 17008
rect 1492 15904 1544 15910
rect 1492 15846 1544 15852
rect 1504 15745 1532 15846
rect 1490 15736 1546 15745
rect 1490 15671 1546 15680
rect 1400 15496 1452 15502
rect 1400 15438 1452 15444
rect 1412 15065 1440 15438
rect 1398 15056 1454 15065
rect 1398 14991 1454 15000
rect 1490 14376 1546 14385
rect 1490 14311 1546 14320
rect 1504 14278 1532 14311
rect 1492 14272 1544 14278
rect 1492 14214 1544 14220
rect 1492 12640 1544 12646
rect 1492 12582 1544 12588
rect 1504 12345 1532 12582
rect 1490 12336 1546 12345
rect 1490 12271 1546 12280
rect 1400 11688 1452 11694
rect 1398 11656 1400 11665
rect 1452 11656 1454 11665
rect 1398 11591 1454 11600
rect 1412 11354 1440 11591
rect 1400 11348 1452 11354
rect 1400 11290 1452 11296
rect 1596 10810 1624 18226
rect 1872 18222 1900 32778
rect 2320 32768 2372 32774
rect 2320 32710 2372 32716
rect 2136 30592 2188 30598
rect 2136 30534 2188 30540
rect 1952 30116 2004 30122
rect 1952 30058 2004 30064
rect 1964 30025 1992 30058
rect 1950 30016 2006 30025
rect 1950 29951 2006 29960
rect 1964 29850 1992 29951
rect 1952 29844 2004 29850
rect 1952 29786 2004 29792
rect 1952 29028 2004 29034
rect 1952 28970 2004 28976
rect 1964 20618 1992 28970
rect 2044 24812 2096 24818
rect 2044 24754 2096 24760
rect 2056 24614 2084 24754
rect 2044 24608 2096 24614
rect 2044 24550 2096 24556
rect 2056 20806 2084 24550
rect 2044 20800 2096 20806
rect 2044 20742 2096 20748
rect 1964 20590 2084 20618
rect 2056 18630 2084 20590
rect 2148 18902 2176 30534
rect 2228 27872 2280 27878
rect 2228 27814 2280 27820
rect 2240 22506 2268 27814
rect 2228 22500 2280 22506
rect 2228 22442 2280 22448
rect 2136 18896 2188 18902
rect 2136 18838 2188 18844
rect 2136 18760 2188 18766
rect 2136 18702 2188 18708
rect 1952 18624 2004 18630
rect 1952 18566 2004 18572
rect 2044 18624 2096 18630
rect 2044 18566 2096 18572
rect 1860 18216 1912 18222
rect 1860 18158 1912 18164
rect 1860 18080 1912 18086
rect 1860 18022 1912 18028
rect 1676 13252 1728 13258
rect 1676 13194 1728 13200
rect 1688 13025 1716 13194
rect 1674 13016 1730 13025
rect 1674 12951 1730 12960
rect 1584 10804 1636 10810
rect 1584 10746 1636 10752
rect 1400 10668 1452 10674
rect 1400 10610 1452 10616
rect 1412 10305 1440 10610
rect 1398 10296 1454 10305
rect 1398 10231 1454 10240
rect 1490 8936 1546 8945
rect 1490 8871 1546 8880
rect 1504 8838 1532 8871
rect 1492 8832 1544 8838
rect 1492 8774 1544 8780
rect 1492 7744 1544 7750
rect 1492 7686 1544 7692
rect 1504 7585 1532 7686
rect 1490 7576 1546 7585
rect 1490 7511 1546 7520
rect 1492 7200 1544 7206
rect 1492 7142 1544 7148
rect 1504 6905 1532 7142
rect 1490 6896 1546 6905
rect 1490 6831 1546 6840
rect 1490 6216 1546 6225
rect 1490 6151 1492 6160
rect 1544 6151 1546 6160
rect 1492 6122 1544 6128
rect 1492 5024 1544 5030
rect 1492 4966 1544 4972
rect 1504 4865 1532 4966
rect 1490 4856 1546 4865
rect 1490 4791 1546 4800
rect 1400 4480 1452 4486
rect 1400 4422 1452 4428
rect 1412 4146 1440 4422
rect 1400 4140 1452 4146
rect 1400 4082 1452 4088
rect 20 3664 72 3670
rect 20 3606 72 3612
rect 32 800 60 3606
rect 664 3392 716 3398
rect 664 3334 716 3340
rect 676 800 704 3334
rect 1412 2825 1440 4082
rect 1872 3534 1900 18022
rect 1964 17678 1992 18566
rect 2148 18465 2176 18702
rect 2332 18698 2360 32710
rect 2412 29504 2464 29510
rect 2412 29446 2464 29452
rect 2320 18692 2372 18698
rect 2320 18634 2372 18640
rect 2134 18456 2190 18465
rect 2134 18391 2190 18400
rect 2424 18154 2452 29446
rect 2412 18148 2464 18154
rect 2412 18090 2464 18096
rect 2608 17882 2636 33254
rect 2780 32904 2832 32910
rect 2780 32846 2832 32852
rect 2792 31958 2820 32846
rect 2884 32570 2912 34711
rect 2872 32564 2924 32570
rect 2872 32506 2924 32512
rect 2976 32026 3004 35391
rect 3238 35200 3294 36000
rect 3882 35200 3938 36000
rect 4526 35306 4582 36000
rect 5170 35306 5226 36000
rect 5814 35306 5870 36000
rect 6458 35306 6514 36000
rect 7746 35306 7802 36000
rect 8390 35306 8446 36000
rect 9034 35306 9090 36000
rect 9678 35306 9734 36000
rect 10322 35306 10378 36000
rect 10966 35306 11022 36000
rect 4526 35278 4660 35306
rect 4526 35200 4582 35278
rect 3896 33658 3924 35200
rect 3884 33652 3936 33658
rect 3884 33594 3936 33600
rect 4632 33522 4660 35278
rect 5170 35278 5488 35306
rect 5170 35200 5226 35278
rect 5460 33538 5488 35278
rect 5814 35278 6040 35306
rect 5814 35200 5870 35278
rect 5460 33522 5580 33538
rect 3976 33516 4028 33522
rect 3976 33458 4028 33464
rect 4620 33516 4672 33522
rect 5460 33516 5592 33522
rect 5460 33510 5540 33516
rect 4620 33458 4672 33464
rect 5540 33458 5592 33464
rect 3056 33448 3108 33454
rect 3056 33390 3108 33396
rect 2964 32020 3016 32026
rect 2964 31962 3016 31968
rect 2780 31952 2832 31958
rect 2780 31894 2832 31900
rect 2964 31816 3016 31822
rect 2964 31758 3016 31764
rect 2976 26450 3004 31758
rect 2964 26444 3016 26450
rect 2964 26386 3016 26392
rect 3068 18358 3096 33390
rect 3988 33318 4016 33458
rect 3976 33312 4028 33318
rect 3976 33254 4028 33260
rect 4632 33114 4660 33458
rect 5552 33114 5580 33458
rect 6012 33114 6040 35278
rect 6458 35278 6776 35306
rect 6458 35200 6514 35278
rect 6748 33658 6776 35278
rect 7746 35278 7972 35306
rect 7746 35200 7802 35278
rect 6736 33652 6788 33658
rect 6736 33594 6788 33600
rect 7944 33522 7972 35278
rect 8390 35278 8524 35306
rect 8390 35200 8446 35278
rect 8496 33522 8524 35278
rect 9034 35278 9352 35306
rect 9034 35200 9090 35278
rect 6368 33516 6420 33522
rect 6368 33458 6420 33464
rect 7932 33516 7984 33522
rect 7932 33458 7984 33464
rect 8484 33516 8536 33522
rect 8484 33458 8536 33464
rect 4620 33108 4672 33114
rect 4620 33050 4672 33056
rect 5540 33108 5592 33114
rect 5540 33050 5592 33056
rect 6000 33108 6052 33114
rect 6000 33050 6052 33056
rect 3516 32904 3568 32910
rect 3516 32846 3568 32852
rect 3424 26512 3476 26518
rect 3424 26454 3476 26460
rect 3436 18358 3464 26454
rect 3528 18426 3556 32846
rect 6092 25152 6144 25158
rect 6092 25094 6144 25100
rect 4068 23724 4120 23730
rect 4068 23666 4120 23672
rect 4080 18426 4108 23666
rect 6104 22642 6132 25094
rect 6092 22636 6144 22642
rect 6092 22578 6144 22584
rect 3516 18420 3568 18426
rect 3516 18362 3568 18368
rect 4068 18420 4120 18426
rect 4068 18362 4120 18368
rect 6380 18358 6408 33458
rect 8024 33312 8076 33318
rect 8024 33254 8076 33260
rect 6582 33212 6890 33232
rect 6582 33210 6588 33212
rect 6644 33210 6668 33212
rect 6724 33210 6748 33212
rect 6804 33210 6828 33212
rect 6884 33210 6890 33212
rect 6644 33158 6646 33210
rect 6826 33158 6828 33210
rect 6582 33156 6588 33158
rect 6644 33156 6668 33158
rect 6724 33156 6748 33158
rect 6804 33156 6828 33158
rect 6884 33156 6890 33158
rect 6582 33136 6890 33156
rect 6460 32768 6512 32774
rect 6460 32710 6512 32716
rect 6472 27470 6500 32710
rect 6582 32124 6890 32144
rect 6582 32122 6588 32124
rect 6644 32122 6668 32124
rect 6724 32122 6748 32124
rect 6804 32122 6828 32124
rect 6884 32122 6890 32124
rect 6644 32070 6646 32122
rect 6826 32070 6828 32122
rect 6582 32068 6588 32070
rect 6644 32068 6668 32070
rect 6724 32068 6748 32070
rect 6804 32068 6828 32070
rect 6884 32068 6890 32070
rect 6582 32048 6890 32068
rect 6582 31036 6890 31056
rect 6582 31034 6588 31036
rect 6644 31034 6668 31036
rect 6724 31034 6748 31036
rect 6804 31034 6828 31036
rect 6884 31034 6890 31036
rect 6644 30982 6646 31034
rect 6826 30982 6828 31034
rect 6582 30980 6588 30982
rect 6644 30980 6668 30982
rect 6724 30980 6748 30982
rect 6804 30980 6828 30982
rect 6884 30980 6890 30982
rect 6582 30960 6890 30980
rect 6582 29948 6890 29968
rect 6582 29946 6588 29948
rect 6644 29946 6668 29948
rect 6724 29946 6748 29948
rect 6804 29946 6828 29948
rect 6884 29946 6890 29948
rect 6644 29894 6646 29946
rect 6826 29894 6828 29946
rect 6582 29892 6588 29894
rect 6644 29892 6668 29894
rect 6724 29892 6748 29894
rect 6804 29892 6828 29894
rect 6884 29892 6890 29894
rect 6582 29872 6890 29892
rect 6582 28860 6890 28880
rect 6582 28858 6588 28860
rect 6644 28858 6668 28860
rect 6724 28858 6748 28860
rect 6804 28858 6828 28860
rect 6884 28858 6890 28860
rect 6644 28806 6646 28858
rect 6826 28806 6828 28858
rect 6582 28804 6588 28806
rect 6644 28804 6668 28806
rect 6724 28804 6748 28806
rect 6804 28804 6828 28806
rect 6884 28804 6890 28806
rect 6582 28784 6890 28804
rect 6582 27772 6890 27792
rect 6582 27770 6588 27772
rect 6644 27770 6668 27772
rect 6724 27770 6748 27772
rect 6804 27770 6828 27772
rect 6884 27770 6890 27772
rect 6644 27718 6646 27770
rect 6826 27718 6828 27770
rect 6582 27716 6588 27718
rect 6644 27716 6668 27718
rect 6724 27716 6748 27718
rect 6804 27716 6828 27718
rect 6884 27716 6890 27718
rect 6582 27696 6890 27716
rect 6460 27464 6512 27470
rect 6460 27406 6512 27412
rect 6582 26684 6890 26704
rect 6582 26682 6588 26684
rect 6644 26682 6668 26684
rect 6724 26682 6748 26684
rect 6804 26682 6828 26684
rect 6884 26682 6890 26684
rect 6644 26630 6646 26682
rect 6826 26630 6828 26682
rect 6582 26628 6588 26630
rect 6644 26628 6668 26630
rect 6724 26628 6748 26630
rect 6804 26628 6828 26630
rect 6884 26628 6890 26630
rect 6582 26608 6890 26628
rect 6582 25596 6890 25616
rect 6582 25594 6588 25596
rect 6644 25594 6668 25596
rect 6724 25594 6748 25596
rect 6804 25594 6828 25596
rect 6884 25594 6890 25596
rect 6644 25542 6646 25594
rect 6826 25542 6828 25594
rect 6582 25540 6588 25542
rect 6644 25540 6668 25542
rect 6724 25540 6748 25542
rect 6804 25540 6828 25542
rect 6884 25540 6890 25542
rect 6582 25520 6890 25540
rect 6582 24508 6890 24528
rect 6582 24506 6588 24508
rect 6644 24506 6668 24508
rect 6724 24506 6748 24508
rect 6804 24506 6828 24508
rect 6884 24506 6890 24508
rect 6644 24454 6646 24506
rect 6826 24454 6828 24506
rect 6582 24452 6588 24454
rect 6644 24452 6668 24454
rect 6724 24452 6748 24454
rect 6804 24452 6828 24454
rect 6884 24452 6890 24454
rect 6582 24432 6890 24452
rect 6582 23420 6890 23440
rect 6582 23418 6588 23420
rect 6644 23418 6668 23420
rect 6724 23418 6748 23420
rect 6804 23418 6828 23420
rect 6884 23418 6890 23420
rect 6644 23366 6646 23418
rect 6826 23366 6828 23418
rect 6582 23364 6588 23366
rect 6644 23364 6668 23366
rect 6724 23364 6748 23366
rect 6804 23364 6828 23366
rect 6884 23364 6890 23366
rect 6582 23344 6890 23364
rect 6582 22332 6890 22352
rect 6582 22330 6588 22332
rect 6644 22330 6668 22332
rect 6724 22330 6748 22332
rect 6804 22330 6828 22332
rect 6884 22330 6890 22332
rect 6644 22278 6646 22330
rect 6826 22278 6828 22330
rect 6582 22276 6588 22278
rect 6644 22276 6668 22278
rect 6724 22276 6748 22278
rect 6804 22276 6828 22278
rect 6884 22276 6890 22278
rect 6582 22256 6890 22276
rect 6582 21244 6890 21264
rect 6582 21242 6588 21244
rect 6644 21242 6668 21244
rect 6724 21242 6748 21244
rect 6804 21242 6828 21244
rect 6884 21242 6890 21244
rect 6644 21190 6646 21242
rect 6826 21190 6828 21242
rect 6582 21188 6588 21190
rect 6644 21188 6668 21190
rect 6724 21188 6748 21190
rect 6804 21188 6828 21190
rect 6884 21188 6890 21190
rect 6582 21168 6890 21188
rect 6582 20156 6890 20176
rect 6582 20154 6588 20156
rect 6644 20154 6668 20156
rect 6724 20154 6748 20156
rect 6804 20154 6828 20156
rect 6884 20154 6890 20156
rect 6644 20102 6646 20154
rect 6826 20102 6828 20154
rect 6582 20100 6588 20102
rect 6644 20100 6668 20102
rect 6724 20100 6748 20102
rect 6804 20100 6828 20102
rect 6884 20100 6890 20102
rect 6582 20080 6890 20100
rect 6582 19068 6890 19088
rect 6582 19066 6588 19068
rect 6644 19066 6668 19068
rect 6724 19066 6748 19068
rect 6804 19066 6828 19068
rect 6884 19066 6890 19068
rect 6644 19014 6646 19066
rect 6826 19014 6828 19066
rect 6582 19012 6588 19014
rect 6644 19012 6668 19014
rect 6724 19012 6748 19014
rect 6804 19012 6828 19014
rect 6884 19012 6890 19014
rect 6582 18992 6890 19012
rect 3056 18352 3108 18358
rect 3056 18294 3108 18300
rect 3424 18352 3476 18358
rect 3424 18294 3476 18300
rect 6368 18352 6420 18358
rect 6368 18294 6420 18300
rect 6920 18352 6972 18358
rect 6920 18294 6972 18300
rect 3608 18284 3660 18290
rect 3608 18226 3660 18232
rect 6460 18284 6512 18290
rect 6460 18226 6512 18232
rect 2964 18080 3016 18086
rect 2964 18022 3016 18028
rect 2596 17876 2648 17882
rect 2596 17818 2648 17824
rect 1952 17672 2004 17678
rect 1952 17614 2004 17620
rect 2504 17604 2556 17610
rect 2504 17546 2556 17552
rect 2412 17536 2464 17542
rect 2412 17478 2464 17484
rect 2044 12844 2096 12850
rect 2044 12786 2096 12792
rect 2056 12646 2084 12786
rect 2044 12640 2096 12646
rect 2044 12582 2096 12588
rect 2056 9382 2084 12582
rect 2044 9376 2096 9382
rect 2044 9318 2096 9324
rect 2044 7404 2096 7410
rect 2044 7346 2096 7352
rect 2056 7206 2084 7346
rect 2044 7200 2096 7206
rect 2044 7142 2096 7148
rect 2056 4486 2084 7142
rect 2044 4480 2096 4486
rect 2044 4422 2096 4428
rect 2044 3936 2096 3942
rect 2044 3878 2096 3884
rect 2056 3534 2084 3878
rect 1860 3528 1912 3534
rect 1860 3470 1912 3476
rect 2044 3528 2096 3534
rect 2044 3470 2096 3476
rect 2424 3058 2452 17478
rect 2516 15706 2544 17546
rect 2504 15700 2556 15706
rect 2504 15642 2556 15648
rect 2976 6322 3004 18022
rect 2964 6316 3016 6322
rect 2964 6258 3016 6264
rect 3056 4140 3108 4146
rect 3056 4082 3108 4088
rect 3068 3942 3096 4082
rect 3056 3936 3108 3942
rect 3056 3878 3108 3884
rect 2964 3392 3016 3398
rect 2964 3334 3016 3340
rect 2412 3052 2464 3058
rect 2412 2994 2464 3000
rect 2976 2990 3004 3334
rect 2964 2984 3016 2990
rect 2964 2926 3016 2932
rect 2596 2916 2648 2922
rect 2596 2858 2648 2864
rect 1952 2848 2004 2854
rect 1398 2816 1454 2825
rect 1952 2790 2004 2796
rect 1398 2751 1454 2760
rect 1400 2508 1452 2514
rect 1400 2450 1452 2456
rect 1412 2394 1440 2450
rect 1320 2366 1440 2394
rect 1320 800 1348 2366
rect 1964 800 1992 2790
rect 2608 2514 2636 2858
rect 2872 2848 2924 2854
rect 2872 2790 2924 2796
rect 2596 2508 2648 2514
rect 2596 2450 2648 2456
rect 2504 2440 2556 2446
rect 2504 2382 2556 2388
rect 2516 2106 2544 2382
rect 2884 2378 2912 2790
rect 2872 2372 2924 2378
rect 2872 2314 2924 2320
rect 2780 2304 2832 2310
rect 2608 2264 2780 2292
rect 2504 2100 2556 2106
rect 2504 2042 2556 2048
rect 2608 800 2636 2264
rect 2780 2246 2832 2252
rect 2884 2145 2912 2314
rect 2870 2136 2926 2145
rect 2870 2071 2926 2080
rect 2976 1465 3004 2926
rect 2962 1456 3018 1465
rect 2962 1391 3018 1400
rect 18 0 74 800
rect 662 0 718 800
rect 1306 0 1362 800
rect 1950 0 2006 800
rect 2594 0 2650 800
rect 2962 776 3018 785
rect 3068 762 3096 3878
rect 3620 2514 3648 18226
rect 6472 6914 6500 18226
rect 6932 18154 6960 18294
rect 7288 18284 7340 18290
rect 7288 18226 7340 18232
rect 6920 18148 6972 18154
rect 6920 18090 6972 18096
rect 6582 17980 6890 18000
rect 6582 17978 6588 17980
rect 6644 17978 6668 17980
rect 6724 17978 6748 17980
rect 6804 17978 6828 17980
rect 6884 17978 6890 17980
rect 6644 17926 6646 17978
rect 6826 17926 6828 17978
rect 6582 17924 6588 17926
rect 6644 17924 6668 17926
rect 6724 17924 6748 17926
rect 6804 17924 6828 17926
rect 6884 17924 6890 17926
rect 6582 17904 6890 17924
rect 6582 16892 6890 16912
rect 6582 16890 6588 16892
rect 6644 16890 6668 16892
rect 6724 16890 6748 16892
rect 6804 16890 6828 16892
rect 6884 16890 6890 16892
rect 6644 16838 6646 16890
rect 6826 16838 6828 16890
rect 6582 16836 6588 16838
rect 6644 16836 6668 16838
rect 6724 16836 6748 16838
rect 6804 16836 6828 16838
rect 6884 16836 6890 16838
rect 6582 16816 6890 16836
rect 6582 15804 6890 15824
rect 6582 15802 6588 15804
rect 6644 15802 6668 15804
rect 6724 15802 6748 15804
rect 6804 15802 6828 15804
rect 6884 15802 6890 15804
rect 6644 15750 6646 15802
rect 6826 15750 6828 15802
rect 6582 15748 6588 15750
rect 6644 15748 6668 15750
rect 6724 15748 6748 15750
rect 6804 15748 6828 15750
rect 6884 15748 6890 15750
rect 6582 15728 6890 15748
rect 6582 14716 6890 14736
rect 6582 14714 6588 14716
rect 6644 14714 6668 14716
rect 6724 14714 6748 14716
rect 6804 14714 6828 14716
rect 6884 14714 6890 14716
rect 6644 14662 6646 14714
rect 6826 14662 6828 14714
rect 6582 14660 6588 14662
rect 6644 14660 6668 14662
rect 6724 14660 6748 14662
rect 6804 14660 6828 14662
rect 6884 14660 6890 14662
rect 6582 14640 6890 14660
rect 6582 13628 6890 13648
rect 6582 13626 6588 13628
rect 6644 13626 6668 13628
rect 6724 13626 6748 13628
rect 6804 13626 6828 13628
rect 6884 13626 6890 13628
rect 6644 13574 6646 13626
rect 6826 13574 6828 13626
rect 6582 13572 6588 13574
rect 6644 13572 6668 13574
rect 6724 13572 6748 13574
rect 6804 13572 6828 13574
rect 6884 13572 6890 13574
rect 6582 13552 6890 13572
rect 6582 12540 6890 12560
rect 6582 12538 6588 12540
rect 6644 12538 6668 12540
rect 6724 12538 6748 12540
rect 6804 12538 6828 12540
rect 6884 12538 6890 12540
rect 6644 12486 6646 12538
rect 6826 12486 6828 12538
rect 6582 12484 6588 12486
rect 6644 12484 6668 12486
rect 6724 12484 6748 12486
rect 6804 12484 6828 12486
rect 6884 12484 6890 12486
rect 6582 12464 6890 12484
rect 6582 11452 6890 11472
rect 6582 11450 6588 11452
rect 6644 11450 6668 11452
rect 6724 11450 6748 11452
rect 6804 11450 6828 11452
rect 6884 11450 6890 11452
rect 6644 11398 6646 11450
rect 6826 11398 6828 11450
rect 6582 11396 6588 11398
rect 6644 11396 6668 11398
rect 6724 11396 6748 11398
rect 6804 11396 6828 11398
rect 6884 11396 6890 11398
rect 6582 11376 6890 11396
rect 6582 10364 6890 10384
rect 6582 10362 6588 10364
rect 6644 10362 6668 10364
rect 6724 10362 6748 10364
rect 6804 10362 6828 10364
rect 6884 10362 6890 10364
rect 6644 10310 6646 10362
rect 6826 10310 6828 10362
rect 6582 10308 6588 10310
rect 6644 10308 6668 10310
rect 6724 10308 6748 10310
rect 6804 10308 6828 10310
rect 6884 10308 6890 10310
rect 6582 10288 6890 10308
rect 6582 9276 6890 9296
rect 6582 9274 6588 9276
rect 6644 9274 6668 9276
rect 6724 9274 6748 9276
rect 6804 9274 6828 9276
rect 6884 9274 6890 9276
rect 6644 9222 6646 9274
rect 6826 9222 6828 9274
rect 6582 9220 6588 9222
rect 6644 9220 6668 9222
rect 6724 9220 6748 9222
rect 6804 9220 6828 9222
rect 6884 9220 6890 9222
rect 6582 9200 6890 9220
rect 6582 8188 6890 8208
rect 6582 8186 6588 8188
rect 6644 8186 6668 8188
rect 6724 8186 6748 8188
rect 6804 8186 6828 8188
rect 6884 8186 6890 8188
rect 6644 8134 6646 8186
rect 6826 8134 6828 8186
rect 6582 8132 6588 8134
rect 6644 8132 6668 8134
rect 6724 8132 6748 8134
rect 6804 8132 6828 8134
rect 6884 8132 6890 8134
rect 6582 8112 6890 8132
rect 6582 7100 6890 7120
rect 6582 7098 6588 7100
rect 6644 7098 6668 7100
rect 6724 7098 6748 7100
rect 6804 7098 6828 7100
rect 6884 7098 6890 7100
rect 6644 7046 6646 7098
rect 6826 7046 6828 7098
rect 6582 7044 6588 7046
rect 6644 7044 6668 7046
rect 6724 7044 6748 7046
rect 6804 7044 6828 7046
rect 6884 7044 6890 7046
rect 6582 7024 6890 7044
rect 6380 6886 6500 6914
rect 4436 3596 4488 3602
rect 4436 3538 4488 3544
rect 4252 3460 4304 3466
rect 4252 3402 4304 3408
rect 3792 3392 3844 3398
rect 3792 3334 3844 3340
rect 4160 3392 4212 3398
rect 4160 3334 4212 3340
rect 3608 2508 3660 2514
rect 3608 2450 3660 2456
rect 3804 2446 3832 3334
rect 3884 2848 3936 2854
rect 3884 2790 3936 2796
rect 3240 2440 3292 2446
rect 3240 2382 3292 2388
rect 3424 2440 3476 2446
rect 3424 2382 3476 2388
rect 3792 2440 3844 2446
rect 3792 2382 3844 2388
rect 3252 2038 3280 2382
rect 3240 2032 3292 2038
rect 3240 1974 3292 1980
rect 3436 1850 3464 2382
rect 3252 1822 3464 1850
rect 3252 800 3280 1822
rect 3896 800 3924 2790
rect 4172 2582 4200 3334
rect 4264 3058 4292 3402
rect 4448 3126 4476 3538
rect 4436 3120 4488 3126
rect 4436 3062 4488 3068
rect 4252 3052 4304 3058
rect 4252 2994 4304 3000
rect 4528 2848 4580 2854
rect 4528 2790 4580 2796
rect 5816 2848 5868 2854
rect 5816 2790 5868 2796
rect 4160 2576 4212 2582
rect 4160 2518 4212 2524
rect 4540 2446 4568 2790
rect 5828 2446 5856 2790
rect 6380 2582 6408 6886
rect 6582 6012 6890 6032
rect 6582 6010 6588 6012
rect 6644 6010 6668 6012
rect 6724 6010 6748 6012
rect 6804 6010 6828 6012
rect 6884 6010 6890 6012
rect 6644 5958 6646 6010
rect 6826 5958 6828 6010
rect 6582 5956 6588 5958
rect 6644 5956 6668 5958
rect 6724 5956 6748 5958
rect 6804 5956 6828 5958
rect 6884 5956 6890 5958
rect 6582 5936 6890 5956
rect 6582 4924 6890 4944
rect 6582 4922 6588 4924
rect 6644 4922 6668 4924
rect 6724 4922 6748 4924
rect 6804 4922 6828 4924
rect 6884 4922 6890 4924
rect 6644 4870 6646 4922
rect 6826 4870 6828 4922
rect 6582 4868 6588 4870
rect 6644 4868 6668 4870
rect 6724 4868 6748 4870
rect 6804 4868 6828 4870
rect 6884 4868 6890 4870
rect 6582 4848 6890 4868
rect 6582 3836 6890 3856
rect 6582 3834 6588 3836
rect 6644 3834 6668 3836
rect 6724 3834 6748 3836
rect 6804 3834 6828 3836
rect 6884 3834 6890 3836
rect 6644 3782 6646 3834
rect 6826 3782 6828 3834
rect 6582 3780 6588 3782
rect 6644 3780 6668 3782
rect 6724 3780 6748 3782
rect 6804 3780 6828 3782
rect 6884 3780 6890 3782
rect 6582 3760 6890 3780
rect 6828 3664 6880 3670
rect 6828 3606 6880 3612
rect 6840 3058 6868 3606
rect 6828 3052 6880 3058
rect 6828 2994 6880 3000
rect 6460 2848 6512 2854
rect 6460 2790 6512 2796
rect 6368 2576 6420 2582
rect 6368 2518 6420 2524
rect 4528 2440 4580 2446
rect 4528 2382 4580 2388
rect 5816 2440 5868 2446
rect 5816 2382 5868 2388
rect 4540 800 4568 2382
rect 5828 800 5856 2382
rect 6472 800 6500 2790
rect 6582 2748 6890 2768
rect 6582 2746 6588 2748
rect 6644 2746 6668 2748
rect 6724 2746 6748 2748
rect 6804 2746 6828 2748
rect 6884 2746 6890 2748
rect 6644 2694 6646 2746
rect 6826 2694 6828 2746
rect 6582 2692 6588 2694
rect 6644 2692 6668 2694
rect 6724 2692 6748 2694
rect 6804 2692 6828 2694
rect 6884 2692 6890 2694
rect 6582 2672 6890 2692
rect 7300 2514 7328 18226
rect 8036 17610 8064 33254
rect 8496 33114 8524 33458
rect 8484 33108 8536 33114
rect 8484 33050 8536 33056
rect 9324 32910 9352 35278
rect 9678 35278 9904 35306
rect 9678 35200 9734 35278
rect 9876 33658 9904 35278
rect 10322 35278 10640 35306
rect 10322 35200 10378 35278
rect 10508 33924 10560 33930
rect 10508 33866 10560 33872
rect 9864 33652 9916 33658
rect 9864 33594 9916 33600
rect 10520 33454 10548 33866
rect 10612 33454 10640 35278
rect 10796 35278 11022 35306
rect 10508 33448 10560 33454
rect 10508 33390 10560 33396
rect 10600 33448 10652 33454
rect 10600 33390 10652 33396
rect 10796 33114 10824 35278
rect 10966 35200 11022 35278
rect 11610 35306 11666 36000
rect 11610 35278 11744 35306
rect 11610 35200 11666 35278
rect 11612 33992 11664 33998
rect 11612 33934 11664 33940
rect 11152 33448 11204 33454
rect 11152 33390 11204 33396
rect 11164 33114 11192 33390
rect 11624 33386 11652 33934
rect 11716 33522 11744 35278
rect 12898 35200 12954 36000
rect 13542 35306 13598 36000
rect 14186 35306 14242 36000
rect 14830 35306 14886 36000
rect 13542 35278 13768 35306
rect 13542 35200 13598 35278
rect 12214 33756 12522 33776
rect 12214 33754 12220 33756
rect 12276 33754 12300 33756
rect 12356 33754 12380 33756
rect 12436 33754 12460 33756
rect 12516 33754 12522 33756
rect 12276 33702 12278 33754
rect 12458 33702 12460 33754
rect 12214 33700 12220 33702
rect 12276 33700 12300 33702
rect 12356 33700 12380 33702
rect 12436 33700 12460 33702
rect 12516 33700 12522 33702
rect 12214 33680 12522 33700
rect 11704 33516 11756 33522
rect 11704 33458 11756 33464
rect 13740 33402 13768 35278
rect 14186 35278 14504 35306
rect 14186 35200 14242 35278
rect 14372 33856 14424 33862
rect 14372 33798 14424 33804
rect 14384 33522 14412 33798
rect 14476 33522 14504 35278
rect 14660 35278 14886 35306
rect 14372 33516 14424 33522
rect 14372 33458 14424 33464
rect 14464 33516 14516 33522
rect 14464 33458 14516 33464
rect 13740 33386 13860 33402
rect 11612 33380 11664 33386
rect 13740 33380 13872 33386
rect 13740 33374 13820 33380
rect 11612 33322 11664 33328
rect 13820 33322 13872 33328
rect 11888 33312 11940 33318
rect 11888 33254 11940 33260
rect 10784 33108 10836 33114
rect 10784 33050 10836 33056
rect 11152 33108 11204 33114
rect 11152 33050 11204 33056
rect 10796 32910 10824 33050
rect 9312 32904 9364 32910
rect 9312 32846 9364 32852
rect 10784 32904 10836 32910
rect 10784 32846 10836 32852
rect 9128 32768 9180 32774
rect 9128 32710 9180 32716
rect 11244 32768 11296 32774
rect 11244 32710 11296 32716
rect 9140 25294 9168 32710
rect 11256 32434 11284 32710
rect 11244 32428 11296 32434
rect 11244 32370 11296 32376
rect 11900 31414 11928 33254
rect 14660 33114 14688 35278
rect 14830 35200 14886 35278
rect 15474 35200 15530 36000
rect 16118 35306 16174 36000
rect 16118 35278 16436 35306
rect 16118 35200 16174 35278
rect 15016 33924 15068 33930
rect 15016 33866 15068 33872
rect 14740 33584 14792 33590
rect 14740 33526 14792 33532
rect 14648 33108 14700 33114
rect 14648 33050 14700 33056
rect 14752 33046 14780 33526
rect 14740 33040 14792 33046
rect 14740 32982 14792 32988
rect 15028 32978 15056 33866
rect 15488 33590 15516 35200
rect 15476 33584 15528 33590
rect 15476 33526 15528 33532
rect 15568 33312 15620 33318
rect 15568 33254 15620 33260
rect 15580 32994 15608 33254
rect 16408 33114 16436 35278
rect 16762 35200 16818 36000
rect 18050 35200 18106 36000
rect 18694 35200 18750 36000
rect 19338 35306 19394 36000
rect 19338 35278 19472 35306
rect 19338 35200 19394 35278
rect 16672 33924 16724 33930
rect 16672 33866 16724 33872
rect 16684 33658 16712 33866
rect 16776 33658 16804 35200
rect 18064 33658 18092 35200
rect 18420 33992 18472 33998
rect 18420 33934 18472 33940
rect 16672 33652 16724 33658
rect 16672 33594 16724 33600
rect 16764 33652 16816 33658
rect 16764 33594 16816 33600
rect 18052 33652 18104 33658
rect 18052 33594 18104 33600
rect 17132 33516 17184 33522
rect 17132 33458 17184 33464
rect 17144 33114 17172 33458
rect 17408 33448 17460 33454
rect 17408 33390 17460 33396
rect 16396 33108 16448 33114
rect 16396 33050 16448 33056
rect 17132 33108 17184 33114
rect 17132 33050 17184 33056
rect 15016 32972 15068 32978
rect 15580 32966 16252 32994
rect 15016 32914 15068 32920
rect 15200 32904 15252 32910
rect 15200 32846 15252 32852
rect 15568 32904 15620 32910
rect 15568 32846 15620 32852
rect 12214 32668 12522 32688
rect 12214 32666 12220 32668
rect 12276 32666 12300 32668
rect 12356 32666 12380 32668
rect 12436 32666 12460 32668
rect 12516 32666 12522 32668
rect 12276 32614 12278 32666
rect 12458 32614 12460 32666
rect 12214 32612 12220 32614
rect 12276 32612 12300 32614
rect 12356 32612 12380 32614
rect 12436 32612 12460 32614
rect 12516 32612 12522 32614
rect 12214 32592 12522 32612
rect 12214 31580 12522 31600
rect 12214 31578 12220 31580
rect 12276 31578 12300 31580
rect 12356 31578 12380 31580
rect 12436 31578 12460 31580
rect 12516 31578 12522 31580
rect 12276 31526 12278 31578
rect 12458 31526 12460 31578
rect 12214 31524 12220 31526
rect 12276 31524 12300 31526
rect 12356 31524 12380 31526
rect 12436 31524 12460 31526
rect 12516 31524 12522 31526
rect 12214 31504 12522 31524
rect 11888 31408 11940 31414
rect 11888 31350 11940 31356
rect 12214 30492 12522 30512
rect 12214 30490 12220 30492
rect 12276 30490 12300 30492
rect 12356 30490 12380 30492
rect 12436 30490 12460 30492
rect 12516 30490 12522 30492
rect 12276 30438 12278 30490
rect 12458 30438 12460 30490
rect 12214 30436 12220 30438
rect 12276 30436 12300 30438
rect 12356 30436 12380 30438
rect 12436 30436 12460 30438
rect 12516 30436 12522 30438
rect 12214 30416 12522 30436
rect 12214 29404 12522 29424
rect 12214 29402 12220 29404
rect 12276 29402 12300 29404
rect 12356 29402 12380 29404
rect 12436 29402 12460 29404
rect 12516 29402 12522 29404
rect 12276 29350 12278 29402
rect 12458 29350 12460 29402
rect 12214 29348 12220 29350
rect 12276 29348 12300 29350
rect 12356 29348 12380 29350
rect 12436 29348 12460 29350
rect 12516 29348 12522 29350
rect 12214 29328 12522 29348
rect 12214 28316 12522 28336
rect 12214 28314 12220 28316
rect 12276 28314 12300 28316
rect 12356 28314 12380 28316
rect 12436 28314 12460 28316
rect 12516 28314 12522 28316
rect 12276 28262 12278 28314
rect 12458 28262 12460 28314
rect 12214 28260 12220 28262
rect 12276 28260 12300 28262
rect 12356 28260 12380 28262
rect 12436 28260 12460 28262
rect 12516 28260 12522 28262
rect 12214 28240 12522 28260
rect 12214 27228 12522 27248
rect 12214 27226 12220 27228
rect 12276 27226 12300 27228
rect 12356 27226 12380 27228
rect 12436 27226 12460 27228
rect 12516 27226 12522 27228
rect 12276 27174 12278 27226
rect 12458 27174 12460 27226
rect 12214 27172 12220 27174
rect 12276 27172 12300 27174
rect 12356 27172 12380 27174
rect 12436 27172 12460 27174
rect 12516 27172 12522 27174
rect 12214 27152 12522 27172
rect 12214 26140 12522 26160
rect 12214 26138 12220 26140
rect 12276 26138 12300 26140
rect 12356 26138 12380 26140
rect 12436 26138 12460 26140
rect 12516 26138 12522 26140
rect 12276 26086 12278 26138
rect 12458 26086 12460 26138
rect 12214 26084 12220 26086
rect 12276 26084 12300 26086
rect 12356 26084 12380 26086
rect 12436 26084 12460 26086
rect 12516 26084 12522 26086
rect 12214 26064 12522 26084
rect 9128 25288 9180 25294
rect 9128 25230 9180 25236
rect 12214 25052 12522 25072
rect 12214 25050 12220 25052
rect 12276 25050 12300 25052
rect 12356 25050 12380 25052
rect 12436 25050 12460 25052
rect 12516 25050 12522 25052
rect 12276 24998 12278 25050
rect 12458 24998 12460 25050
rect 12214 24996 12220 24998
rect 12276 24996 12300 24998
rect 12356 24996 12380 24998
rect 12436 24996 12460 24998
rect 12516 24996 12522 24998
rect 12214 24976 12522 24996
rect 12214 23964 12522 23984
rect 12214 23962 12220 23964
rect 12276 23962 12300 23964
rect 12356 23962 12380 23964
rect 12436 23962 12460 23964
rect 12516 23962 12522 23964
rect 12276 23910 12278 23962
rect 12458 23910 12460 23962
rect 12214 23908 12220 23910
rect 12276 23908 12300 23910
rect 12356 23908 12380 23910
rect 12436 23908 12460 23910
rect 12516 23908 12522 23910
rect 12214 23888 12522 23908
rect 12214 22876 12522 22896
rect 12214 22874 12220 22876
rect 12276 22874 12300 22876
rect 12356 22874 12380 22876
rect 12436 22874 12460 22876
rect 12516 22874 12522 22876
rect 12276 22822 12278 22874
rect 12458 22822 12460 22874
rect 12214 22820 12220 22822
rect 12276 22820 12300 22822
rect 12356 22820 12380 22822
rect 12436 22820 12460 22822
rect 12516 22820 12522 22822
rect 12214 22800 12522 22820
rect 12214 21788 12522 21808
rect 12214 21786 12220 21788
rect 12276 21786 12300 21788
rect 12356 21786 12380 21788
rect 12436 21786 12460 21788
rect 12516 21786 12522 21788
rect 12276 21734 12278 21786
rect 12458 21734 12460 21786
rect 12214 21732 12220 21734
rect 12276 21732 12300 21734
rect 12356 21732 12380 21734
rect 12436 21732 12460 21734
rect 12516 21732 12522 21734
rect 12214 21712 12522 21732
rect 12214 20700 12522 20720
rect 12214 20698 12220 20700
rect 12276 20698 12300 20700
rect 12356 20698 12380 20700
rect 12436 20698 12460 20700
rect 12516 20698 12522 20700
rect 12276 20646 12278 20698
rect 12458 20646 12460 20698
rect 12214 20644 12220 20646
rect 12276 20644 12300 20646
rect 12356 20644 12380 20646
rect 12436 20644 12460 20646
rect 12516 20644 12522 20646
rect 12214 20624 12522 20644
rect 12214 19612 12522 19632
rect 12214 19610 12220 19612
rect 12276 19610 12300 19612
rect 12356 19610 12380 19612
rect 12436 19610 12460 19612
rect 12516 19610 12522 19612
rect 12276 19558 12278 19610
rect 12458 19558 12460 19610
rect 12214 19556 12220 19558
rect 12276 19556 12300 19558
rect 12356 19556 12380 19558
rect 12436 19556 12460 19558
rect 12516 19556 12522 19558
rect 12214 19536 12522 19556
rect 12900 18828 12952 18834
rect 12900 18770 12952 18776
rect 12214 18524 12522 18544
rect 12214 18522 12220 18524
rect 12276 18522 12300 18524
rect 12356 18522 12380 18524
rect 12436 18522 12460 18524
rect 12516 18522 12522 18524
rect 12276 18470 12278 18522
rect 12458 18470 12460 18522
rect 12214 18468 12220 18470
rect 12276 18468 12300 18470
rect 12356 18468 12380 18470
rect 12436 18468 12460 18470
rect 12516 18468 12522 18470
rect 12214 18448 12522 18468
rect 12912 18426 12940 18770
rect 12900 18420 12952 18426
rect 12900 18362 12952 18368
rect 8116 18352 8168 18358
rect 8116 18294 8168 18300
rect 8024 17604 8076 17610
rect 8024 17546 8076 17552
rect 8128 3738 8156 18294
rect 15212 18290 15240 32846
rect 15292 32836 15344 32842
rect 15292 32778 15344 32784
rect 15304 31929 15332 32778
rect 15580 32570 15608 32846
rect 15568 32564 15620 32570
rect 15568 32506 15620 32512
rect 15290 31920 15346 31929
rect 15290 31855 15346 31864
rect 16224 18426 16252 32966
rect 16580 26852 16632 26858
rect 16580 26794 16632 26800
rect 16592 24138 16620 26794
rect 16580 24132 16632 24138
rect 16580 24074 16632 24080
rect 17224 19168 17276 19174
rect 17224 19110 17276 19116
rect 17236 18766 17264 19110
rect 17224 18760 17276 18766
rect 17224 18702 17276 18708
rect 16212 18420 16264 18426
rect 16212 18362 16264 18368
rect 15200 18284 15252 18290
rect 15200 18226 15252 18232
rect 15844 18284 15896 18290
rect 15844 18226 15896 18232
rect 16764 18284 16816 18290
rect 16764 18226 16816 18232
rect 17040 18284 17092 18290
rect 17040 18226 17092 18232
rect 15856 17882 15884 18226
rect 16776 18086 16804 18226
rect 16948 18148 17000 18154
rect 16948 18090 17000 18096
rect 16764 18080 16816 18086
rect 16764 18022 16816 18028
rect 16776 17882 16804 18022
rect 15844 17876 15896 17882
rect 15844 17818 15896 17824
rect 16764 17876 16816 17882
rect 16764 17818 16816 17824
rect 16856 17876 16908 17882
rect 16856 17818 16908 17824
rect 12214 17436 12522 17456
rect 12214 17434 12220 17436
rect 12276 17434 12300 17436
rect 12356 17434 12380 17436
rect 12436 17434 12460 17436
rect 12516 17434 12522 17436
rect 12276 17382 12278 17434
rect 12458 17382 12460 17434
rect 12214 17380 12220 17382
rect 12276 17380 12300 17382
rect 12356 17380 12380 17382
rect 12436 17380 12460 17382
rect 12516 17380 12522 17382
rect 12214 17360 12522 17380
rect 12214 16348 12522 16368
rect 12214 16346 12220 16348
rect 12276 16346 12300 16348
rect 12356 16346 12380 16348
rect 12436 16346 12460 16348
rect 12516 16346 12522 16348
rect 12276 16294 12278 16346
rect 12458 16294 12460 16346
rect 12214 16292 12220 16294
rect 12276 16292 12300 16294
rect 12356 16292 12380 16294
rect 12436 16292 12460 16294
rect 12516 16292 12522 16294
rect 12214 16272 12522 16292
rect 12214 15260 12522 15280
rect 12214 15258 12220 15260
rect 12276 15258 12300 15260
rect 12356 15258 12380 15260
rect 12436 15258 12460 15260
rect 12516 15258 12522 15260
rect 12276 15206 12278 15258
rect 12458 15206 12460 15258
rect 12214 15204 12220 15206
rect 12276 15204 12300 15206
rect 12356 15204 12380 15206
rect 12436 15204 12460 15206
rect 12516 15204 12522 15206
rect 12214 15184 12522 15204
rect 11704 14884 11756 14890
rect 11704 14826 11756 14832
rect 11716 14414 11744 14826
rect 11704 14408 11756 14414
rect 11704 14350 11756 14356
rect 12214 14172 12522 14192
rect 12214 14170 12220 14172
rect 12276 14170 12300 14172
rect 12356 14170 12380 14172
rect 12436 14170 12460 14172
rect 12516 14170 12522 14172
rect 12276 14118 12278 14170
rect 12458 14118 12460 14170
rect 12214 14116 12220 14118
rect 12276 14116 12300 14118
rect 12356 14116 12380 14118
rect 12436 14116 12460 14118
rect 12516 14116 12522 14118
rect 12214 14096 12522 14116
rect 12214 13084 12522 13104
rect 12214 13082 12220 13084
rect 12276 13082 12300 13084
rect 12356 13082 12380 13084
rect 12436 13082 12460 13084
rect 12516 13082 12522 13084
rect 12276 13030 12278 13082
rect 12458 13030 12460 13082
rect 12214 13028 12220 13030
rect 12276 13028 12300 13030
rect 12356 13028 12380 13030
rect 12436 13028 12460 13030
rect 12516 13028 12522 13030
rect 12214 13008 12522 13028
rect 12214 11996 12522 12016
rect 12214 11994 12220 11996
rect 12276 11994 12300 11996
rect 12356 11994 12380 11996
rect 12436 11994 12460 11996
rect 12516 11994 12522 11996
rect 12276 11942 12278 11994
rect 12458 11942 12460 11994
rect 12214 11940 12220 11942
rect 12276 11940 12300 11942
rect 12356 11940 12380 11942
rect 12436 11940 12460 11942
rect 12516 11940 12522 11942
rect 12214 11920 12522 11940
rect 12214 10908 12522 10928
rect 12214 10906 12220 10908
rect 12276 10906 12300 10908
rect 12356 10906 12380 10908
rect 12436 10906 12460 10908
rect 12516 10906 12522 10908
rect 12276 10854 12278 10906
rect 12458 10854 12460 10906
rect 12214 10852 12220 10854
rect 12276 10852 12300 10854
rect 12356 10852 12380 10854
rect 12436 10852 12460 10854
rect 12516 10852 12522 10854
rect 12214 10832 12522 10852
rect 12214 9820 12522 9840
rect 12214 9818 12220 9820
rect 12276 9818 12300 9820
rect 12356 9818 12380 9820
rect 12436 9818 12460 9820
rect 12516 9818 12522 9820
rect 12276 9766 12278 9818
rect 12458 9766 12460 9818
rect 12214 9764 12220 9766
rect 12276 9764 12300 9766
rect 12356 9764 12380 9766
rect 12436 9764 12460 9766
rect 12516 9764 12522 9766
rect 12214 9744 12522 9764
rect 12214 8732 12522 8752
rect 12214 8730 12220 8732
rect 12276 8730 12300 8732
rect 12356 8730 12380 8732
rect 12436 8730 12460 8732
rect 12516 8730 12522 8732
rect 12276 8678 12278 8730
rect 12458 8678 12460 8730
rect 12214 8676 12220 8678
rect 12276 8676 12300 8678
rect 12356 8676 12380 8678
rect 12436 8676 12460 8678
rect 12516 8676 12522 8678
rect 12214 8656 12522 8676
rect 10968 7880 11020 7886
rect 10968 7822 11020 7828
rect 10980 5370 11008 7822
rect 12214 7644 12522 7664
rect 12214 7642 12220 7644
rect 12276 7642 12300 7644
rect 12356 7642 12380 7644
rect 12436 7642 12460 7644
rect 12516 7642 12522 7644
rect 12276 7590 12278 7642
rect 12458 7590 12460 7642
rect 12214 7588 12220 7590
rect 12276 7588 12300 7590
rect 12356 7588 12380 7590
rect 12436 7588 12460 7590
rect 12516 7588 12522 7590
rect 12214 7568 12522 7588
rect 12214 6556 12522 6576
rect 12214 6554 12220 6556
rect 12276 6554 12300 6556
rect 12356 6554 12380 6556
rect 12436 6554 12460 6556
rect 12516 6554 12522 6556
rect 12276 6502 12278 6554
rect 12458 6502 12460 6554
rect 12214 6500 12220 6502
rect 12276 6500 12300 6502
rect 12356 6500 12380 6502
rect 12436 6500 12460 6502
rect 12516 6500 12522 6502
rect 12214 6480 12522 6500
rect 12214 5468 12522 5488
rect 12214 5466 12220 5468
rect 12276 5466 12300 5468
rect 12356 5466 12380 5468
rect 12436 5466 12460 5468
rect 12516 5466 12522 5468
rect 12276 5414 12278 5466
rect 12458 5414 12460 5466
rect 12214 5412 12220 5414
rect 12276 5412 12300 5414
rect 12356 5412 12380 5414
rect 12436 5412 12460 5414
rect 12516 5412 12522 5414
rect 12214 5392 12522 5412
rect 10968 5364 11020 5370
rect 10968 5306 11020 5312
rect 13636 5228 13688 5234
rect 13636 5170 13688 5176
rect 12214 4380 12522 4400
rect 12214 4378 12220 4380
rect 12276 4378 12300 4380
rect 12356 4378 12380 4380
rect 12436 4378 12460 4380
rect 12516 4378 12522 4380
rect 12276 4326 12278 4378
rect 12458 4326 12460 4378
rect 12214 4324 12220 4326
rect 12276 4324 12300 4326
rect 12356 4324 12380 4326
rect 12436 4324 12460 4326
rect 12516 4324 12522 4326
rect 12214 4304 12522 4324
rect 11612 4004 11664 4010
rect 11612 3946 11664 3952
rect 8116 3732 8168 3738
rect 8116 3674 8168 3680
rect 7748 3052 7800 3058
rect 7748 2994 7800 3000
rect 7288 2508 7340 2514
rect 7288 2450 7340 2456
rect 7104 2304 7156 2310
rect 7104 2246 7156 2252
rect 7116 800 7144 2246
rect 7760 800 7788 2994
rect 8128 2446 8156 3674
rect 11624 3058 11652 3946
rect 11704 3392 11756 3398
rect 11704 3334 11756 3340
rect 11612 3052 11664 3058
rect 11612 2994 11664 3000
rect 11716 2990 11744 3334
rect 12214 3292 12522 3312
rect 12214 3290 12220 3292
rect 12276 3290 12300 3292
rect 12356 3290 12380 3292
rect 12436 3290 12460 3292
rect 12516 3290 12522 3292
rect 12276 3238 12278 3290
rect 12458 3238 12460 3290
rect 12214 3236 12220 3238
rect 12276 3236 12300 3238
rect 12356 3236 12380 3238
rect 12436 3236 12460 3238
rect 12516 3236 12522 3238
rect 12214 3216 12522 3236
rect 13648 3194 13676 5170
rect 14556 3732 14608 3738
rect 14556 3674 14608 3680
rect 13728 3664 13780 3670
rect 13728 3606 13780 3612
rect 13740 3194 13768 3606
rect 13636 3188 13688 3194
rect 13636 3130 13688 3136
rect 13728 3188 13780 3194
rect 13728 3130 13780 3136
rect 13544 3052 13596 3058
rect 13544 2994 13596 3000
rect 14372 3052 14424 3058
rect 14372 2994 14424 3000
rect 11704 2984 11756 2990
rect 11704 2926 11756 2932
rect 10232 2916 10284 2922
rect 10232 2858 10284 2864
rect 10968 2916 11020 2922
rect 10968 2858 11020 2864
rect 12440 2916 12492 2922
rect 12440 2858 12492 2864
rect 9036 2848 9088 2854
rect 9036 2790 9088 2796
rect 9048 2446 9076 2790
rect 10244 2446 10272 2858
rect 10980 2446 11008 2858
rect 12452 2446 12480 2858
rect 13556 2854 13584 2994
rect 12992 2848 13044 2854
rect 12992 2790 13044 2796
rect 13544 2848 13596 2854
rect 13544 2790 13596 2796
rect 13728 2848 13780 2854
rect 13728 2790 13780 2796
rect 13004 2514 13032 2790
rect 12992 2508 13044 2514
rect 12992 2450 13044 2456
rect 8024 2440 8076 2446
rect 8024 2382 8076 2388
rect 8116 2440 8168 2446
rect 8116 2382 8168 2388
rect 9036 2440 9088 2446
rect 9036 2382 9088 2388
rect 10232 2440 10284 2446
rect 10232 2382 10284 2388
rect 10968 2440 11020 2446
rect 10968 2382 11020 2388
rect 12440 2440 12492 2446
rect 12440 2382 12492 2388
rect 8036 1834 8064 2382
rect 8392 2304 8444 2310
rect 8392 2246 8444 2252
rect 8024 1828 8076 1834
rect 8024 1770 8076 1776
rect 8404 800 8432 2246
rect 9048 800 9076 2382
rect 9680 2304 9732 2310
rect 9680 2246 9732 2252
rect 9692 800 9720 2246
rect 10980 800 11008 2382
rect 11888 2372 11940 2378
rect 11888 2314 11940 2320
rect 11152 2304 11204 2310
rect 11152 2246 11204 2252
rect 11612 2304 11664 2310
rect 11612 2246 11664 2252
rect 11164 1970 11192 2246
rect 11152 1964 11204 1970
rect 11152 1906 11204 1912
rect 11624 800 11652 2246
rect 11900 2106 11928 2314
rect 12072 2304 12124 2310
rect 12072 2246 12124 2252
rect 12900 2304 12952 2310
rect 12900 2246 12952 2252
rect 11888 2100 11940 2106
rect 11888 2042 11940 2048
rect 12084 1170 12112 2246
rect 12214 2204 12522 2224
rect 12214 2202 12220 2204
rect 12276 2202 12300 2204
rect 12356 2202 12380 2204
rect 12436 2202 12460 2204
rect 12516 2202 12522 2204
rect 12276 2150 12278 2202
rect 12458 2150 12460 2202
rect 12214 2148 12220 2150
rect 12276 2148 12300 2150
rect 12356 2148 12380 2150
rect 12436 2148 12460 2150
rect 12516 2148 12522 2150
rect 12214 2128 12522 2148
rect 12084 1142 12296 1170
rect 12268 800 12296 1142
rect 12912 800 12940 2246
rect 13556 800 13584 2790
rect 13740 2446 13768 2790
rect 14384 2650 14412 2994
rect 14372 2644 14424 2650
rect 14372 2586 14424 2592
rect 14568 2582 14596 3674
rect 16672 3528 16724 3534
rect 16672 3470 16724 3476
rect 15200 2848 15252 2854
rect 15200 2790 15252 2796
rect 14556 2576 14608 2582
rect 14556 2518 14608 2524
rect 13728 2440 13780 2446
rect 13728 2382 13780 2388
rect 14832 2440 14884 2446
rect 14832 2382 14884 2388
rect 13740 2310 13768 2382
rect 13728 2304 13780 2310
rect 13728 2246 13780 2252
rect 14188 2304 14240 2310
rect 14188 2246 14240 2252
rect 14200 800 14228 2246
rect 14844 800 14872 2382
rect 15212 1834 15240 2790
rect 16120 2304 16172 2310
rect 16120 2246 16172 2252
rect 15200 1828 15252 1834
rect 15200 1770 15252 1776
rect 16132 800 16160 2246
rect 16684 2038 16712 3470
rect 16764 2440 16816 2446
rect 16764 2382 16816 2388
rect 16672 2032 16724 2038
rect 16672 1974 16724 1980
rect 16776 800 16804 2382
rect 16868 2378 16896 17818
rect 16960 2446 16988 18090
rect 17052 17882 17080 18226
rect 17040 17876 17092 17882
rect 17040 17818 17092 17824
rect 17420 17678 17448 33390
rect 17776 33380 17828 33386
rect 17776 33322 17828 33328
rect 17788 25974 17816 33322
rect 17846 33212 18154 33232
rect 17846 33210 17852 33212
rect 17908 33210 17932 33212
rect 17988 33210 18012 33212
rect 18068 33210 18092 33212
rect 18148 33210 18154 33212
rect 17908 33158 17910 33210
rect 18090 33158 18092 33210
rect 17846 33156 17852 33158
rect 17908 33156 17932 33158
rect 17988 33156 18012 33158
rect 18068 33156 18092 33158
rect 18148 33156 18154 33158
rect 17846 33136 18154 33156
rect 17846 32124 18154 32144
rect 17846 32122 17852 32124
rect 17908 32122 17932 32124
rect 17988 32122 18012 32124
rect 18068 32122 18092 32124
rect 18148 32122 18154 32124
rect 17908 32070 17910 32122
rect 18090 32070 18092 32122
rect 17846 32068 17852 32070
rect 17908 32068 17932 32070
rect 17988 32068 18012 32070
rect 18068 32068 18092 32070
rect 18148 32068 18154 32070
rect 17846 32048 18154 32068
rect 17846 31036 18154 31056
rect 17846 31034 17852 31036
rect 17908 31034 17932 31036
rect 17988 31034 18012 31036
rect 18068 31034 18092 31036
rect 18148 31034 18154 31036
rect 17908 30982 17910 31034
rect 18090 30982 18092 31034
rect 17846 30980 17852 30982
rect 17908 30980 17932 30982
rect 17988 30980 18012 30982
rect 18068 30980 18092 30982
rect 18148 30980 18154 30982
rect 17846 30960 18154 30980
rect 17846 29948 18154 29968
rect 17846 29946 17852 29948
rect 17908 29946 17932 29948
rect 17988 29946 18012 29948
rect 18068 29946 18092 29948
rect 18148 29946 18154 29948
rect 17908 29894 17910 29946
rect 18090 29894 18092 29946
rect 17846 29892 17852 29894
rect 17908 29892 17932 29894
rect 17988 29892 18012 29894
rect 18068 29892 18092 29894
rect 18148 29892 18154 29894
rect 17846 29872 18154 29892
rect 17846 28860 18154 28880
rect 17846 28858 17852 28860
rect 17908 28858 17932 28860
rect 17988 28858 18012 28860
rect 18068 28858 18092 28860
rect 18148 28858 18154 28860
rect 17908 28806 17910 28858
rect 18090 28806 18092 28858
rect 17846 28804 17852 28806
rect 17908 28804 17932 28806
rect 17988 28804 18012 28806
rect 18068 28804 18092 28806
rect 18148 28804 18154 28806
rect 17846 28784 18154 28804
rect 17846 27772 18154 27792
rect 17846 27770 17852 27772
rect 17908 27770 17932 27772
rect 17988 27770 18012 27772
rect 18068 27770 18092 27772
rect 18148 27770 18154 27772
rect 17908 27718 17910 27770
rect 18090 27718 18092 27770
rect 17846 27716 17852 27718
rect 17908 27716 17932 27718
rect 17988 27716 18012 27718
rect 18068 27716 18092 27718
rect 18148 27716 18154 27718
rect 17846 27696 18154 27716
rect 18432 27334 18460 33934
rect 18604 33584 18656 33590
rect 18604 33526 18656 33532
rect 18512 33312 18564 33318
rect 18512 33254 18564 33260
rect 18524 32842 18552 33254
rect 18512 32836 18564 32842
rect 18512 32778 18564 32784
rect 18512 32428 18564 32434
rect 18512 32370 18564 32376
rect 18524 30190 18552 32370
rect 18512 30184 18564 30190
rect 18512 30126 18564 30132
rect 18420 27328 18472 27334
rect 18420 27270 18472 27276
rect 18432 27130 18460 27270
rect 18420 27124 18472 27130
rect 18420 27066 18472 27072
rect 18236 26988 18288 26994
rect 18236 26930 18288 26936
rect 17846 26684 18154 26704
rect 17846 26682 17852 26684
rect 17908 26682 17932 26684
rect 17988 26682 18012 26684
rect 18068 26682 18092 26684
rect 18148 26682 18154 26684
rect 17908 26630 17910 26682
rect 18090 26630 18092 26682
rect 17846 26628 17852 26630
rect 17908 26628 17932 26630
rect 17988 26628 18012 26630
rect 18068 26628 18092 26630
rect 18148 26628 18154 26630
rect 17846 26608 18154 26628
rect 18248 26586 18276 26930
rect 18236 26580 18288 26586
rect 18236 26522 18288 26528
rect 17776 25968 17828 25974
rect 17776 25910 17828 25916
rect 18420 25696 18472 25702
rect 18420 25638 18472 25644
rect 17846 25596 18154 25616
rect 17846 25594 17852 25596
rect 17908 25594 17932 25596
rect 17988 25594 18012 25596
rect 18068 25594 18092 25596
rect 18148 25594 18154 25596
rect 17908 25542 17910 25594
rect 18090 25542 18092 25594
rect 17846 25540 17852 25542
rect 17908 25540 17932 25542
rect 17988 25540 18012 25542
rect 18068 25540 18092 25542
rect 18148 25540 18154 25542
rect 17846 25520 18154 25540
rect 18432 25430 18460 25638
rect 18420 25424 18472 25430
rect 18420 25366 18472 25372
rect 17846 24508 18154 24528
rect 17846 24506 17852 24508
rect 17908 24506 17932 24508
rect 17988 24506 18012 24508
rect 18068 24506 18092 24508
rect 18148 24506 18154 24508
rect 17908 24454 17910 24506
rect 18090 24454 18092 24506
rect 17846 24452 17852 24454
rect 17908 24452 17932 24454
rect 17988 24452 18012 24454
rect 18068 24452 18092 24454
rect 18148 24452 18154 24454
rect 17846 24432 18154 24452
rect 17846 23420 18154 23440
rect 17846 23418 17852 23420
rect 17908 23418 17932 23420
rect 17988 23418 18012 23420
rect 18068 23418 18092 23420
rect 18148 23418 18154 23420
rect 17908 23366 17910 23418
rect 18090 23366 18092 23418
rect 17846 23364 17852 23366
rect 17908 23364 17932 23366
rect 17988 23364 18012 23366
rect 18068 23364 18092 23366
rect 18148 23364 18154 23366
rect 17846 23344 18154 23364
rect 17846 22332 18154 22352
rect 17846 22330 17852 22332
rect 17908 22330 17932 22332
rect 17988 22330 18012 22332
rect 18068 22330 18092 22332
rect 18148 22330 18154 22332
rect 17908 22278 17910 22330
rect 18090 22278 18092 22330
rect 17846 22276 17852 22278
rect 17908 22276 17932 22278
rect 17988 22276 18012 22278
rect 18068 22276 18092 22278
rect 18148 22276 18154 22278
rect 17846 22256 18154 22276
rect 18616 22094 18644 33526
rect 18708 33114 18736 35200
rect 18972 33856 19024 33862
rect 18972 33798 19024 33804
rect 18788 33516 18840 33522
rect 18788 33458 18840 33464
rect 18696 33108 18748 33114
rect 18696 33050 18748 33056
rect 18800 31754 18828 33458
rect 18800 31726 18920 31754
rect 18696 26784 18748 26790
rect 18696 26726 18748 26732
rect 18708 26382 18736 26726
rect 18696 26376 18748 26382
rect 18696 26318 18748 26324
rect 18708 25906 18736 26318
rect 18696 25900 18748 25906
rect 18696 25842 18748 25848
rect 18616 22066 18828 22094
rect 17846 21244 18154 21264
rect 17846 21242 17852 21244
rect 17908 21242 17932 21244
rect 17988 21242 18012 21244
rect 18068 21242 18092 21244
rect 18148 21242 18154 21244
rect 17908 21190 17910 21242
rect 18090 21190 18092 21242
rect 17846 21188 17852 21190
rect 17908 21188 17932 21190
rect 17988 21188 18012 21190
rect 18068 21188 18092 21190
rect 18148 21188 18154 21190
rect 17846 21168 18154 21188
rect 17846 20156 18154 20176
rect 17846 20154 17852 20156
rect 17908 20154 17932 20156
rect 17988 20154 18012 20156
rect 18068 20154 18092 20156
rect 18148 20154 18154 20156
rect 17908 20102 17910 20154
rect 18090 20102 18092 20154
rect 17846 20100 17852 20102
rect 17908 20100 17932 20102
rect 17988 20100 18012 20102
rect 18068 20100 18092 20102
rect 18148 20100 18154 20102
rect 17846 20080 18154 20100
rect 17960 19780 18012 19786
rect 17960 19722 18012 19728
rect 17972 19446 18000 19722
rect 17960 19440 18012 19446
rect 17960 19382 18012 19388
rect 18328 19372 18380 19378
rect 18328 19314 18380 19320
rect 17846 19068 18154 19088
rect 17846 19066 17852 19068
rect 17908 19066 17932 19068
rect 17988 19066 18012 19068
rect 18068 19066 18092 19068
rect 18148 19066 18154 19068
rect 17908 19014 17910 19066
rect 18090 19014 18092 19066
rect 17846 19012 17852 19014
rect 17908 19012 17932 19014
rect 17988 19012 18012 19014
rect 18068 19012 18092 19014
rect 18148 19012 18154 19014
rect 17846 18992 18154 19012
rect 18236 18692 18288 18698
rect 18236 18634 18288 18640
rect 17500 18148 17552 18154
rect 17500 18090 17552 18096
rect 17408 17672 17460 17678
rect 17408 17614 17460 17620
rect 17408 17536 17460 17542
rect 17408 17478 17460 17484
rect 17420 17338 17448 17478
rect 17408 17332 17460 17338
rect 17408 17274 17460 17280
rect 17512 16574 17540 18090
rect 17846 17980 18154 18000
rect 17846 17978 17852 17980
rect 17908 17978 17932 17980
rect 17988 17978 18012 17980
rect 18068 17978 18092 17980
rect 18148 17978 18154 17980
rect 17908 17926 17910 17978
rect 18090 17926 18092 17978
rect 17846 17924 17852 17926
rect 17908 17924 17932 17926
rect 17988 17924 18012 17926
rect 18068 17924 18092 17926
rect 18148 17924 18154 17926
rect 17846 17904 18154 17924
rect 17776 17604 17828 17610
rect 17776 17546 17828 17552
rect 17684 17196 17736 17202
rect 17684 17138 17736 17144
rect 17696 16794 17724 17138
rect 17684 16788 17736 16794
rect 17684 16730 17736 16736
rect 17512 16546 17632 16574
rect 17316 9988 17368 9994
rect 17316 9930 17368 9936
rect 17132 3596 17184 3602
rect 17132 3538 17184 3544
rect 17144 3058 17172 3538
rect 17224 3528 17276 3534
rect 17224 3470 17276 3476
rect 17132 3052 17184 3058
rect 17132 2994 17184 3000
rect 16948 2440 17000 2446
rect 16948 2382 17000 2388
rect 16856 2372 16908 2378
rect 16856 2314 16908 2320
rect 17236 2106 17264 3470
rect 17328 2650 17356 9930
rect 17604 4486 17632 16546
rect 17696 13258 17724 16730
rect 17684 13252 17736 13258
rect 17684 13194 17736 13200
rect 17788 12850 17816 17546
rect 17846 16892 18154 16912
rect 17846 16890 17852 16892
rect 17908 16890 17932 16892
rect 17988 16890 18012 16892
rect 18068 16890 18092 16892
rect 18148 16890 18154 16892
rect 17908 16838 17910 16890
rect 18090 16838 18092 16890
rect 17846 16836 17852 16838
rect 17908 16836 17932 16838
rect 17988 16836 18012 16838
rect 18068 16836 18092 16838
rect 18148 16836 18154 16838
rect 17846 16816 18154 16836
rect 17846 15804 18154 15824
rect 17846 15802 17852 15804
rect 17908 15802 17932 15804
rect 17988 15802 18012 15804
rect 18068 15802 18092 15804
rect 18148 15802 18154 15804
rect 17908 15750 17910 15802
rect 18090 15750 18092 15802
rect 17846 15748 17852 15750
rect 17908 15748 17932 15750
rect 17988 15748 18012 15750
rect 18068 15748 18092 15750
rect 18148 15748 18154 15750
rect 17846 15728 18154 15748
rect 17846 14716 18154 14736
rect 17846 14714 17852 14716
rect 17908 14714 17932 14716
rect 17988 14714 18012 14716
rect 18068 14714 18092 14716
rect 18148 14714 18154 14716
rect 17908 14662 17910 14714
rect 18090 14662 18092 14714
rect 17846 14660 17852 14662
rect 17908 14660 17932 14662
rect 17988 14660 18012 14662
rect 18068 14660 18092 14662
rect 18148 14660 18154 14662
rect 17846 14640 18154 14660
rect 17846 13628 18154 13648
rect 17846 13626 17852 13628
rect 17908 13626 17932 13628
rect 17988 13626 18012 13628
rect 18068 13626 18092 13628
rect 18148 13626 18154 13628
rect 17908 13574 17910 13626
rect 18090 13574 18092 13626
rect 17846 13572 17852 13574
rect 17908 13572 17932 13574
rect 17988 13572 18012 13574
rect 18068 13572 18092 13574
rect 18148 13572 18154 13574
rect 17846 13552 18154 13572
rect 17776 12844 17828 12850
rect 17776 12786 17828 12792
rect 17846 12540 18154 12560
rect 17846 12538 17852 12540
rect 17908 12538 17932 12540
rect 17988 12538 18012 12540
rect 18068 12538 18092 12540
rect 18148 12538 18154 12540
rect 17908 12486 17910 12538
rect 18090 12486 18092 12538
rect 17846 12484 17852 12486
rect 17908 12484 17932 12486
rect 17988 12484 18012 12486
rect 18068 12484 18092 12486
rect 18148 12484 18154 12486
rect 17846 12464 18154 12484
rect 17846 11452 18154 11472
rect 17846 11450 17852 11452
rect 17908 11450 17932 11452
rect 17988 11450 18012 11452
rect 18068 11450 18092 11452
rect 18148 11450 18154 11452
rect 17908 11398 17910 11450
rect 18090 11398 18092 11450
rect 17846 11396 17852 11398
rect 17908 11396 17932 11398
rect 17988 11396 18012 11398
rect 18068 11396 18092 11398
rect 18148 11396 18154 11398
rect 17846 11376 18154 11396
rect 17846 10364 18154 10384
rect 17846 10362 17852 10364
rect 17908 10362 17932 10364
rect 17988 10362 18012 10364
rect 18068 10362 18092 10364
rect 18148 10362 18154 10364
rect 17908 10310 17910 10362
rect 18090 10310 18092 10362
rect 17846 10308 17852 10310
rect 17908 10308 17932 10310
rect 17988 10308 18012 10310
rect 18068 10308 18092 10310
rect 18148 10308 18154 10310
rect 17846 10288 18154 10308
rect 17846 9276 18154 9296
rect 17846 9274 17852 9276
rect 17908 9274 17932 9276
rect 17988 9274 18012 9276
rect 18068 9274 18092 9276
rect 18148 9274 18154 9276
rect 17908 9222 17910 9274
rect 18090 9222 18092 9274
rect 17846 9220 17852 9222
rect 17908 9220 17932 9222
rect 17988 9220 18012 9222
rect 18068 9220 18092 9222
rect 18148 9220 18154 9222
rect 17846 9200 18154 9220
rect 18248 8974 18276 18634
rect 18236 8968 18288 8974
rect 18236 8910 18288 8916
rect 17846 8188 18154 8208
rect 17846 8186 17852 8188
rect 17908 8186 17932 8188
rect 17988 8186 18012 8188
rect 18068 8186 18092 8188
rect 18148 8186 18154 8188
rect 17908 8134 17910 8186
rect 18090 8134 18092 8186
rect 17846 8132 17852 8134
rect 17908 8132 17932 8134
rect 17988 8132 18012 8134
rect 18068 8132 18092 8134
rect 18148 8132 18154 8134
rect 17846 8112 18154 8132
rect 17846 7100 18154 7120
rect 17846 7098 17852 7100
rect 17908 7098 17932 7100
rect 17988 7098 18012 7100
rect 18068 7098 18092 7100
rect 18148 7098 18154 7100
rect 17908 7046 17910 7098
rect 18090 7046 18092 7098
rect 17846 7044 17852 7046
rect 17908 7044 17932 7046
rect 17988 7044 18012 7046
rect 18068 7044 18092 7046
rect 18148 7044 18154 7046
rect 17846 7024 18154 7044
rect 18340 6914 18368 19314
rect 18800 18766 18828 22066
rect 18788 18760 18840 18766
rect 18788 18702 18840 18708
rect 18696 18692 18748 18698
rect 18696 18634 18748 18640
rect 18604 17604 18656 17610
rect 18604 17546 18656 17552
rect 18616 17134 18644 17546
rect 18604 17128 18656 17134
rect 18604 17070 18656 17076
rect 18708 16574 18736 18634
rect 18892 17882 18920 31726
rect 18984 18086 19012 33798
rect 19444 33522 19472 35278
rect 19982 35200 20038 36000
rect 20626 35200 20682 36000
rect 21270 35200 21326 36000
rect 21914 35200 21970 36000
rect 23202 35306 23258 36000
rect 23032 35278 23258 35306
rect 20260 33924 20312 33930
rect 20260 33866 20312 33872
rect 19432 33516 19484 33522
rect 19432 33458 19484 33464
rect 19800 33448 19852 33454
rect 19800 33390 19852 33396
rect 19340 33380 19392 33386
rect 19340 33322 19392 33328
rect 19248 32904 19300 32910
rect 19248 32846 19300 32852
rect 19064 26988 19116 26994
rect 19064 26930 19116 26936
rect 19076 26042 19104 26930
rect 19064 26036 19116 26042
rect 19064 25978 19116 25984
rect 19260 25498 19288 32846
rect 19352 32842 19380 33322
rect 19340 32836 19392 32842
rect 19340 32778 19392 32784
rect 19340 27124 19392 27130
rect 19340 27066 19392 27072
rect 19248 25492 19300 25498
rect 19248 25434 19300 25440
rect 19248 19168 19300 19174
rect 19248 19110 19300 19116
rect 19064 18624 19116 18630
rect 19064 18566 19116 18572
rect 18972 18080 19024 18086
rect 18972 18022 19024 18028
rect 18880 17876 18932 17882
rect 18880 17818 18932 17824
rect 19076 16574 19104 18566
rect 18708 16546 18828 16574
rect 18512 16108 18564 16114
rect 18512 16050 18564 16056
rect 18524 15162 18552 16050
rect 18512 15156 18564 15162
rect 18512 15098 18564 15104
rect 18512 9580 18564 9586
rect 18512 9522 18564 9528
rect 18524 9382 18552 9522
rect 18512 9376 18564 9382
rect 18512 9318 18564 9324
rect 18248 6886 18368 6914
rect 17846 6012 18154 6032
rect 17846 6010 17852 6012
rect 17908 6010 17932 6012
rect 17988 6010 18012 6012
rect 18068 6010 18092 6012
rect 18148 6010 18154 6012
rect 17908 5958 17910 6010
rect 18090 5958 18092 6010
rect 17846 5956 17852 5958
rect 17908 5956 17932 5958
rect 17988 5956 18012 5958
rect 18068 5956 18092 5958
rect 18148 5956 18154 5958
rect 17846 5936 18154 5956
rect 17776 5160 17828 5166
rect 17776 5102 17828 5108
rect 17788 4758 17816 5102
rect 17846 4924 18154 4944
rect 17846 4922 17852 4924
rect 17908 4922 17932 4924
rect 17988 4922 18012 4924
rect 18068 4922 18092 4924
rect 18148 4922 18154 4924
rect 17908 4870 17910 4922
rect 18090 4870 18092 4922
rect 17846 4868 17852 4870
rect 17908 4868 17932 4870
rect 17988 4868 18012 4870
rect 18068 4868 18092 4870
rect 18148 4868 18154 4870
rect 17846 4848 18154 4868
rect 17776 4752 17828 4758
rect 17776 4694 17828 4700
rect 17592 4480 17644 4486
rect 17592 4422 17644 4428
rect 17846 3836 18154 3856
rect 17846 3834 17852 3836
rect 17908 3834 17932 3836
rect 17988 3834 18012 3836
rect 18068 3834 18092 3836
rect 18148 3834 18154 3836
rect 17908 3782 17910 3834
rect 18090 3782 18092 3834
rect 17846 3780 17852 3782
rect 17908 3780 17932 3782
rect 17988 3780 18012 3782
rect 18068 3780 18092 3782
rect 18148 3780 18154 3782
rect 17846 3760 18154 3780
rect 17408 3664 17460 3670
rect 17408 3606 17460 3612
rect 17420 3058 17448 3606
rect 17776 3460 17828 3466
rect 17776 3402 17828 3408
rect 17500 3392 17552 3398
rect 17500 3334 17552 3340
rect 17408 3052 17460 3058
rect 17408 2994 17460 3000
rect 17316 2644 17368 2650
rect 17316 2586 17368 2592
rect 17512 2446 17540 3334
rect 17788 3126 17816 3402
rect 17776 3120 17828 3126
rect 17776 3062 17828 3068
rect 17846 2748 18154 2768
rect 17846 2746 17852 2748
rect 17908 2746 17932 2748
rect 17988 2746 18012 2748
rect 18068 2746 18092 2748
rect 18148 2746 18154 2748
rect 17908 2694 17910 2746
rect 18090 2694 18092 2746
rect 17846 2692 17852 2694
rect 17908 2692 17932 2694
rect 17988 2692 18012 2694
rect 18068 2692 18092 2694
rect 18148 2692 18154 2694
rect 17846 2672 18154 2692
rect 17500 2440 17552 2446
rect 17500 2382 17552 2388
rect 18052 2440 18104 2446
rect 18052 2382 18104 2388
rect 17408 2304 17460 2310
rect 17408 2246 17460 2252
rect 17224 2100 17276 2106
rect 17224 2042 17276 2048
rect 17420 800 17448 2246
rect 18064 800 18092 2382
rect 18248 1902 18276 6886
rect 18524 3670 18552 9318
rect 18512 3664 18564 3670
rect 18512 3606 18564 3612
rect 18328 3052 18380 3058
rect 18328 2994 18380 3000
rect 18512 3052 18564 3058
rect 18512 2994 18564 3000
rect 18340 2650 18368 2994
rect 18328 2644 18380 2650
rect 18328 2586 18380 2592
rect 18524 1970 18552 2994
rect 18696 2508 18748 2514
rect 18696 2450 18748 2456
rect 18512 1964 18564 1970
rect 18512 1906 18564 1912
rect 18236 1896 18288 1902
rect 18236 1838 18288 1844
rect 18708 800 18736 2450
rect 18800 2378 18828 16546
rect 18892 16546 19104 16574
rect 18892 11626 18920 16546
rect 18972 15020 19024 15026
rect 18972 14962 19024 14968
rect 18984 14822 19012 14962
rect 18972 14816 19024 14822
rect 18972 14758 19024 14764
rect 18880 11620 18932 11626
rect 18880 11562 18932 11568
rect 18984 8362 19012 14758
rect 19260 11778 19288 19110
rect 19076 11750 19288 11778
rect 18972 8356 19024 8362
rect 18972 8298 19024 8304
rect 19076 3505 19104 11750
rect 19248 11620 19300 11626
rect 19248 11562 19300 11568
rect 19062 3496 19118 3505
rect 19062 3431 19118 3440
rect 19156 3460 19208 3466
rect 19156 3402 19208 3408
rect 18880 3392 18932 3398
rect 18880 3334 18932 3340
rect 18892 2446 18920 3334
rect 19168 2514 19196 3402
rect 19260 2990 19288 11562
rect 19352 8906 19380 27066
rect 19708 26376 19760 26382
rect 19708 26318 19760 26324
rect 19616 25900 19668 25906
rect 19616 25842 19668 25848
rect 19628 25362 19656 25842
rect 19616 25356 19668 25362
rect 19616 25298 19668 25304
rect 19720 25226 19748 26318
rect 19708 25220 19760 25226
rect 19708 25162 19760 25168
rect 19812 22094 19840 33390
rect 20272 28218 20300 33866
rect 20640 33522 20668 35200
rect 21284 33522 21312 35200
rect 23032 33658 23060 35278
rect 23202 35200 23258 35278
rect 23846 35306 23902 36000
rect 24490 35306 24546 36000
rect 25134 35306 25190 36000
rect 25778 35306 25834 36000
rect 26422 35306 26478 36000
rect 27066 35306 27122 36000
rect 28354 35306 28410 36000
rect 23846 35278 23980 35306
rect 23846 35200 23902 35278
rect 23478 33756 23786 33776
rect 23478 33754 23484 33756
rect 23540 33754 23564 33756
rect 23620 33754 23644 33756
rect 23700 33754 23724 33756
rect 23780 33754 23786 33756
rect 23540 33702 23542 33754
rect 23722 33702 23724 33754
rect 23478 33700 23484 33702
rect 23540 33700 23564 33702
rect 23620 33700 23644 33702
rect 23700 33700 23724 33702
rect 23780 33700 23786 33702
rect 23478 33680 23786 33700
rect 23952 33658 23980 35278
rect 24490 35278 24716 35306
rect 24490 35200 24546 35278
rect 23020 33652 23072 33658
rect 23020 33594 23072 33600
rect 23940 33652 23992 33658
rect 23940 33594 23992 33600
rect 20628 33516 20680 33522
rect 20628 33458 20680 33464
rect 21272 33516 21324 33522
rect 21272 33458 21324 33464
rect 20640 33114 20668 33458
rect 24492 33448 24544 33454
rect 24492 33390 24544 33396
rect 21916 33312 21968 33318
rect 21916 33254 21968 33260
rect 20628 33108 20680 33114
rect 20628 33050 20680 33056
rect 21928 32910 21956 33254
rect 21916 32904 21968 32910
rect 21916 32846 21968 32852
rect 23478 32668 23786 32688
rect 23478 32666 23484 32668
rect 23540 32666 23564 32668
rect 23620 32666 23644 32668
rect 23700 32666 23724 32668
rect 23780 32666 23786 32668
rect 23540 32614 23542 32666
rect 23722 32614 23724 32666
rect 23478 32612 23484 32614
rect 23540 32612 23564 32614
rect 23620 32612 23644 32614
rect 23700 32612 23724 32614
rect 23780 32612 23786 32614
rect 23478 32592 23786 32612
rect 23478 31580 23786 31600
rect 23478 31578 23484 31580
rect 23540 31578 23564 31580
rect 23620 31578 23644 31580
rect 23700 31578 23724 31580
rect 23780 31578 23786 31580
rect 23540 31526 23542 31578
rect 23722 31526 23724 31578
rect 23478 31524 23484 31526
rect 23540 31524 23564 31526
rect 23620 31524 23644 31526
rect 23700 31524 23724 31526
rect 23780 31524 23786 31526
rect 23478 31504 23786 31524
rect 22100 31136 22152 31142
rect 22100 31078 22152 31084
rect 22112 30938 22140 31078
rect 22100 30932 22152 30938
rect 22100 30874 22152 30880
rect 23478 30492 23786 30512
rect 23478 30490 23484 30492
rect 23540 30490 23564 30492
rect 23620 30490 23644 30492
rect 23700 30490 23724 30492
rect 23780 30490 23786 30492
rect 23540 30438 23542 30490
rect 23722 30438 23724 30490
rect 23478 30436 23484 30438
rect 23540 30436 23564 30438
rect 23620 30436 23644 30438
rect 23700 30436 23724 30438
rect 23780 30436 23786 30438
rect 23478 30416 23786 30436
rect 23478 29404 23786 29424
rect 23478 29402 23484 29404
rect 23540 29402 23564 29404
rect 23620 29402 23644 29404
rect 23700 29402 23724 29404
rect 23780 29402 23786 29404
rect 23540 29350 23542 29402
rect 23722 29350 23724 29402
rect 23478 29348 23484 29350
rect 23540 29348 23564 29350
rect 23620 29348 23644 29350
rect 23700 29348 23724 29350
rect 23780 29348 23786 29350
rect 23478 29328 23786 29348
rect 23478 28316 23786 28336
rect 23478 28314 23484 28316
rect 23540 28314 23564 28316
rect 23620 28314 23644 28316
rect 23700 28314 23724 28316
rect 23780 28314 23786 28316
rect 23540 28262 23542 28314
rect 23722 28262 23724 28314
rect 23478 28260 23484 28262
rect 23540 28260 23564 28262
rect 23620 28260 23644 28262
rect 23700 28260 23724 28262
rect 23780 28260 23786 28262
rect 23478 28240 23786 28260
rect 20260 28212 20312 28218
rect 20260 28154 20312 28160
rect 19984 27600 20036 27606
rect 19984 27542 20036 27548
rect 19996 26994 20024 27542
rect 20272 27470 20300 28154
rect 20076 27464 20128 27470
rect 20076 27406 20128 27412
rect 20260 27464 20312 27470
rect 20260 27406 20312 27412
rect 20628 27464 20680 27470
rect 20628 27406 20680 27412
rect 20088 27130 20116 27406
rect 20076 27124 20128 27130
rect 20076 27066 20128 27072
rect 20272 26994 20300 27406
rect 19892 26988 19944 26994
rect 19892 26930 19944 26936
rect 19984 26988 20036 26994
rect 19984 26930 20036 26936
rect 20260 26988 20312 26994
rect 20260 26930 20312 26936
rect 19904 26042 19932 26930
rect 19996 26602 20024 26930
rect 20640 26926 20668 27406
rect 21180 27396 21232 27402
rect 21180 27338 21232 27344
rect 20812 27328 20864 27334
rect 20812 27270 20864 27276
rect 20628 26920 20680 26926
rect 20628 26862 20680 26868
rect 20260 26852 20312 26858
rect 20260 26794 20312 26800
rect 19996 26574 20116 26602
rect 20088 26382 20116 26574
rect 20272 26382 20300 26794
rect 20352 26784 20404 26790
rect 20352 26726 20404 26732
rect 20364 26518 20392 26726
rect 20352 26512 20404 26518
rect 20352 26454 20404 26460
rect 20076 26376 20128 26382
rect 20076 26318 20128 26324
rect 20260 26376 20312 26382
rect 20260 26318 20312 26324
rect 19892 26036 19944 26042
rect 19892 25978 19944 25984
rect 19984 25900 20036 25906
rect 19984 25842 20036 25848
rect 19996 25498 20024 25842
rect 20088 25770 20116 26318
rect 20272 25906 20300 26318
rect 20364 26246 20392 26454
rect 20824 26382 20852 27270
rect 21192 26586 21220 27338
rect 21640 27328 21692 27334
rect 21640 27270 21692 27276
rect 21652 27062 21680 27270
rect 23478 27228 23786 27248
rect 23478 27226 23484 27228
rect 23540 27226 23564 27228
rect 23620 27226 23644 27228
rect 23700 27226 23724 27228
rect 23780 27226 23786 27228
rect 23540 27174 23542 27226
rect 23722 27174 23724 27226
rect 23478 27172 23484 27174
rect 23540 27172 23564 27174
rect 23620 27172 23644 27174
rect 23700 27172 23724 27174
rect 23780 27172 23786 27174
rect 23478 27152 23786 27172
rect 21640 27056 21692 27062
rect 21640 26998 21692 27004
rect 21916 26988 21968 26994
rect 21916 26930 21968 26936
rect 21928 26790 21956 26930
rect 21916 26784 21968 26790
rect 21916 26726 21968 26732
rect 21088 26580 21140 26586
rect 21088 26522 21140 26528
rect 21180 26580 21232 26586
rect 21180 26522 21232 26528
rect 21100 26382 21128 26522
rect 21928 26450 21956 26726
rect 21916 26444 21968 26450
rect 21916 26386 21968 26392
rect 20812 26376 20864 26382
rect 20812 26318 20864 26324
rect 21088 26376 21140 26382
rect 21088 26318 21140 26324
rect 20352 26240 20404 26246
rect 20352 26182 20404 26188
rect 20904 26240 20956 26246
rect 20904 26182 20956 26188
rect 21456 26240 21508 26246
rect 21456 26182 21508 26188
rect 20260 25900 20312 25906
rect 20260 25842 20312 25848
rect 20076 25764 20128 25770
rect 20076 25706 20128 25712
rect 19984 25492 20036 25498
rect 19984 25434 20036 25440
rect 20272 24954 20300 25842
rect 20364 25702 20392 26182
rect 20916 25906 20944 26182
rect 20904 25900 20956 25906
rect 20904 25842 20956 25848
rect 20916 25786 20944 25842
rect 21468 25838 21496 26182
rect 23478 26140 23786 26160
rect 23478 26138 23484 26140
rect 23540 26138 23564 26140
rect 23620 26138 23644 26140
rect 23700 26138 23724 26140
rect 23780 26138 23786 26140
rect 23540 26086 23542 26138
rect 23722 26086 23724 26138
rect 23478 26084 23484 26086
rect 23540 26084 23564 26086
rect 23620 26084 23644 26086
rect 23700 26084 23724 26086
rect 23780 26084 23786 26086
rect 23478 26064 23786 26084
rect 20824 25758 20944 25786
rect 21456 25832 21508 25838
rect 21456 25774 21508 25780
rect 20352 25696 20404 25702
rect 20352 25638 20404 25644
rect 20364 25498 20392 25638
rect 20352 25492 20404 25498
rect 20352 25434 20404 25440
rect 20352 25356 20404 25362
rect 20352 25298 20404 25304
rect 20364 25226 20392 25298
rect 20824 25294 20852 25758
rect 20996 25696 21048 25702
rect 20996 25638 21048 25644
rect 20628 25288 20680 25294
rect 20812 25288 20864 25294
rect 20680 25236 20760 25242
rect 20628 25230 20760 25236
rect 20812 25230 20864 25236
rect 20352 25220 20404 25226
rect 20640 25214 20760 25230
rect 20352 25162 20404 25168
rect 20364 25106 20392 25162
rect 20732 25158 20760 25214
rect 20720 25152 20772 25158
rect 20364 25078 20484 25106
rect 20720 25094 20772 25100
rect 20260 24948 20312 24954
rect 20260 24890 20312 24896
rect 20456 24614 20484 25078
rect 20444 24608 20496 24614
rect 20444 24550 20496 24556
rect 20456 24070 20484 24550
rect 20444 24064 20496 24070
rect 20444 24006 20496 24012
rect 19812 22066 19932 22094
rect 19524 18284 19576 18290
rect 19524 18226 19576 18232
rect 19616 18284 19668 18290
rect 19616 18226 19668 18232
rect 19432 17604 19484 17610
rect 19432 17546 19484 17552
rect 19340 8900 19392 8906
rect 19340 8842 19392 8848
rect 19248 2984 19300 2990
rect 19248 2926 19300 2932
rect 19340 2848 19392 2854
rect 19340 2790 19392 2796
rect 19156 2508 19208 2514
rect 19156 2450 19208 2456
rect 18880 2440 18932 2446
rect 18880 2382 18932 2388
rect 18788 2372 18840 2378
rect 18788 2314 18840 2320
rect 19352 800 19380 2790
rect 19444 2582 19472 17546
rect 19432 2576 19484 2582
rect 19432 2518 19484 2524
rect 19536 2514 19564 18226
rect 19628 18154 19656 18226
rect 19616 18148 19668 18154
rect 19616 18090 19668 18096
rect 19904 17270 19932 22066
rect 20732 19446 20760 25094
rect 20824 23594 20852 25230
rect 21008 25158 21036 25638
rect 20996 25152 21048 25158
rect 20996 25094 21048 25100
rect 23478 25052 23786 25072
rect 23478 25050 23484 25052
rect 23540 25050 23564 25052
rect 23620 25050 23644 25052
rect 23700 25050 23724 25052
rect 23780 25050 23786 25052
rect 23540 24998 23542 25050
rect 23722 24998 23724 25050
rect 23478 24996 23484 24998
rect 23540 24996 23564 24998
rect 23620 24996 23644 24998
rect 23700 24996 23724 24998
rect 23780 24996 23786 24998
rect 23478 24976 23786 24996
rect 23478 23964 23786 23984
rect 23478 23962 23484 23964
rect 23540 23962 23564 23964
rect 23620 23962 23644 23964
rect 23700 23962 23724 23964
rect 23780 23962 23786 23964
rect 23540 23910 23542 23962
rect 23722 23910 23724 23962
rect 23478 23908 23484 23910
rect 23540 23908 23564 23910
rect 23620 23908 23644 23910
rect 23700 23908 23724 23910
rect 23780 23908 23786 23910
rect 23478 23888 23786 23908
rect 20812 23588 20864 23594
rect 20812 23530 20864 23536
rect 23478 22876 23786 22896
rect 23478 22874 23484 22876
rect 23540 22874 23564 22876
rect 23620 22874 23644 22876
rect 23700 22874 23724 22876
rect 23780 22874 23786 22876
rect 23540 22822 23542 22874
rect 23722 22822 23724 22874
rect 23478 22820 23484 22822
rect 23540 22820 23564 22822
rect 23620 22820 23644 22822
rect 23700 22820 23724 22822
rect 23780 22820 23786 22822
rect 23478 22800 23786 22820
rect 23478 21788 23786 21808
rect 23478 21786 23484 21788
rect 23540 21786 23564 21788
rect 23620 21786 23644 21788
rect 23700 21786 23724 21788
rect 23780 21786 23786 21788
rect 23540 21734 23542 21786
rect 23722 21734 23724 21786
rect 23478 21732 23484 21734
rect 23540 21732 23564 21734
rect 23620 21732 23644 21734
rect 23700 21732 23724 21734
rect 23780 21732 23786 21734
rect 23478 21712 23786 21732
rect 23478 20700 23786 20720
rect 23478 20698 23484 20700
rect 23540 20698 23564 20700
rect 23620 20698 23644 20700
rect 23700 20698 23724 20700
rect 23780 20698 23786 20700
rect 23540 20646 23542 20698
rect 23722 20646 23724 20698
rect 23478 20644 23484 20646
rect 23540 20644 23564 20646
rect 23620 20644 23644 20646
rect 23700 20644 23724 20646
rect 23780 20644 23786 20646
rect 23478 20624 23786 20644
rect 23478 19612 23786 19632
rect 23478 19610 23484 19612
rect 23540 19610 23564 19612
rect 23620 19610 23644 19612
rect 23700 19610 23724 19612
rect 23780 19610 23786 19612
rect 23540 19558 23542 19610
rect 23722 19558 23724 19610
rect 23478 19556 23484 19558
rect 23540 19556 23564 19558
rect 23620 19556 23644 19558
rect 23700 19556 23724 19558
rect 23780 19556 23786 19558
rect 23478 19536 23786 19556
rect 20720 19440 20772 19446
rect 20720 19382 20772 19388
rect 20732 18766 20760 19382
rect 20720 18760 20772 18766
rect 20720 18702 20772 18708
rect 22100 18692 22152 18698
rect 22100 18634 22152 18640
rect 19984 18624 20036 18630
rect 19984 18566 20036 18572
rect 20812 18624 20864 18630
rect 20812 18566 20864 18572
rect 19996 18358 20024 18566
rect 19984 18352 20036 18358
rect 19984 18294 20036 18300
rect 19892 17264 19944 17270
rect 19892 17206 19944 17212
rect 19996 6118 20024 18294
rect 19984 6112 20036 6118
rect 19984 6054 20036 6060
rect 20352 4548 20404 4554
rect 20352 4490 20404 4496
rect 19708 3460 19760 3466
rect 19708 3402 19760 3408
rect 19720 3194 19748 3402
rect 20364 3194 20392 4490
rect 20536 3732 20588 3738
rect 20536 3674 20588 3680
rect 19708 3188 19760 3194
rect 19708 3130 19760 3136
rect 20352 3188 20404 3194
rect 20352 3130 20404 3136
rect 20548 2514 20576 3674
rect 20824 2922 20852 18566
rect 21824 3052 21876 3058
rect 21824 2994 21876 3000
rect 21916 3052 21968 3058
rect 21916 2994 21968 3000
rect 20812 2916 20864 2922
rect 20812 2858 20864 2864
rect 21836 2650 21864 2994
rect 21824 2644 21876 2650
rect 21824 2586 21876 2592
rect 19524 2508 19576 2514
rect 19524 2450 19576 2456
rect 20536 2508 20588 2514
rect 20536 2450 20588 2456
rect 19984 2304 20036 2310
rect 19984 2246 20036 2252
rect 21272 2304 21324 2310
rect 21272 2246 21324 2252
rect 19996 800 20024 2246
rect 21284 800 21312 2246
rect 21928 800 21956 2994
rect 22112 2446 22140 18634
rect 23478 18524 23786 18544
rect 23478 18522 23484 18524
rect 23540 18522 23564 18524
rect 23620 18522 23644 18524
rect 23700 18522 23724 18524
rect 23780 18522 23786 18524
rect 23540 18470 23542 18522
rect 23722 18470 23724 18522
rect 23478 18468 23484 18470
rect 23540 18468 23564 18470
rect 23620 18468 23644 18470
rect 23700 18468 23724 18470
rect 23780 18468 23786 18470
rect 23478 18448 23786 18468
rect 24504 18358 24532 33390
rect 24688 33114 24716 35278
rect 25134 35278 25452 35306
rect 25134 35200 25190 35278
rect 25424 33114 25452 35278
rect 25778 35278 26096 35306
rect 25778 35200 25834 35278
rect 26068 33658 26096 35278
rect 26422 35278 26556 35306
rect 26422 35200 26478 35278
rect 26528 33658 26556 35278
rect 27066 35278 27292 35306
rect 27066 35200 27122 35278
rect 26056 33652 26108 33658
rect 26056 33594 26108 33600
rect 26516 33652 26568 33658
rect 26516 33594 26568 33600
rect 25872 33516 25924 33522
rect 25872 33458 25924 33464
rect 24676 33108 24728 33114
rect 24676 33050 24728 33056
rect 25412 33108 25464 33114
rect 25412 33050 25464 33056
rect 24860 32564 24912 32570
rect 24860 32506 24912 32512
rect 24872 27130 24900 32506
rect 24860 27124 24912 27130
rect 24860 27066 24912 27072
rect 25136 25832 25188 25838
rect 25136 25774 25188 25780
rect 24492 18352 24544 18358
rect 24492 18294 24544 18300
rect 22836 18080 22888 18086
rect 22836 18022 22888 18028
rect 22848 3194 22876 18022
rect 23478 17436 23786 17456
rect 23478 17434 23484 17436
rect 23540 17434 23564 17436
rect 23620 17434 23644 17436
rect 23700 17434 23724 17436
rect 23780 17434 23786 17436
rect 23540 17382 23542 17434
rect 23722 17382 23724 17434
rect 23478 17380 23484 17382
rect 23540 17380 23564 17382
rect 23620 17380 23644 17382
rect 23700 17380 23724 17382
rect 23780 17380 23786 17382
rect 23478 17360 23786 17380
rect 23478 16348 23786 16368
rect 23478 16346 23484 16348
rect 23540 16346 23564 16348
rect 23620 16346 23644 16348
rect 23700 16346 23724 16348
rect 23780 16346 23786 16348
rect 23540 16294 23542 16346
rect 23722 16294 23724 16346
rect 23478 16292 23484 16294
rect 23540 16292 23564 16294
rect 23620 16292 23644 16294
rect 23700 16292 23724 16294
rect 23780 16292 23786 16294
rect 23478 16272 23786 16292
rect 23478 15260 23786 15280
rect 23478 15258 23484 15260
rect 23540 15258 23564 15260
rect 23620 15258 23644 15260
rect 23700 15258 23724 15260
rect 23780 15258 23786 15260
rect 23540 15206 23542 15258
rect 23722 15206 23724 15258
rect 23478 15204 23484 15206
rect 23540 15204 23564 15206
rect 23620 15204 23644 15206
rect 23700 15204 23724 15206
rect 23780 15204 23786 15206
rect 23478 15184 23786 15204
rect 23478 14172 23786 14192
rect 23478 14170 23484 14172
rect 23540 14170 23564 14172
rect 23620 14170 23644 14172
rect 23700 14170 23724 14172
rect 23780 14170 23786 14172
rect 23540 14118 23542 14170
rect 23722 14118 23724 14170
rect 23478 14116 23484 14118
rect 23540 14116 23564 14118
rect 23620 14116 23644 14118
rect 23700 14116 23724 14118
rect 23780 14116 23786 14118
rect 23478 14096 23786 14116
rect 23478 13084 23786 13104
rect 23478 13082 23484 13084
rect 23540 13082 23564 13084
rect 23620 13082 23644 13084
rect 23700 13082 23724 13084
rect 23780 13082 23786 13084
rect 23540 13030 23542 13082
rect 23722 13030 23724 13082
rect 23478 13028 23484 13030
rect 23540 13028 23564 13030
rect 23620 13028 23644 13030
rect 23700 13028 23724 13030
rect 23780 13028 23786 13030
rect 23478 13008 23786 13028
rect 23478 11996 23786 12016
rect 23478 11994 23484 11996
rect 23540 11994 23564 11996
rect 23620 11994 23644 11996
rect 23700 11994 23724 11996
rect 23780 11994 23786 11996
rect 23540 11942 23542 11994
rect 23722 11942 23724 11994
rect 23478 11940 23484 11942
rect 23540 11940 23564 11942
rect 23620 11940 23644 11942
rect 23700 11940 23724 11942
rect 23780 11940 23786 11942
rect 23478 11920 23786 11940
rect 23478 10908 23786 10928
rect 23478 10906 23484 10908
rect 23540 10906 23564 10908
rect 23620 10906 23644 10908
rect 23700 10906 23724 10908
rect 23780 10906 23786 10908
rect 23540 10854 23542 10906
rect 23722 10854 23724 10906
rect 23478 10852 23484 10854
rect 23540 10852 23564 10854
rect 23620 10852 23644 10854
rect 23700 10852 23724 10854
rect 23780 10852 23786 10854
rect 23478 10832 23786 10852
rect 23478 9820 23786 9840
rect 23478 9818 23484 9820
rect 23540 9818 23564 9820
rect 23620 9818 23644 9820
rect 23700 9818 23724 9820
rect 23780 9818 23786 9820
rect 23540 9766 23542 9818
rect 23722 9766 23724 9818
rect 23478 9764 23484 9766
rect 23540 9764 23564 9766
rect 23620 9764 23644 9766
rect 23700 9764 23724 9766
rect 23780 9764 23786 9766
rect 23478 9744 23786 9764
rect 23478 8732 23786 8752
rect 23478 8730 23484 8732
rect 23540 8730 23564 8732
rect 23620 8730 23644 8732
rect 23700 8730 23724 8732
rect 23780 8730 23786 8732
rect 23540 8678 23542 8730
rect 23722 8678 23724 8730
rect 23478 8676 23484 8678
rect 23540 8676 23564 8678
rect 23620 8676 23644 8678
rect 23700 8676 23724 8678
rect 23780 8676 23786 8678
rect 23478 8656 23786 8676
rect 23478 7644 23786 7664
rect 23478 7642 23484 7644
rect 23540 7642 23564 7644
rect 23620 7642 23644 7644
rect 23700 7642 23724 7644
rect 23780 7642 23786 7644
rect 23540 7590 23542 7642
rect 23722 7590 23724 7642
rect 23478 7588 23484 7590
rect 23540 7588 23564 7590
rect 23620 7588 23644 7590
rect 23700 7588 23724 7590
rect 23780 7588 23786 7590
rect 23478 7568 23786 7588
rect 23478 6556 23786 6576
rect 23478 6554 23484 6556
rect 23540 6554 23564 6556
rect 23620 6554 23644 6556
rect 23700 6554 23724 6556
rect 23780 6554 23786 6556
rect 23540 6502 23542 6554
rect 23722 6502 23724 6554
rect 23478 6500 23484 6502
rect 23540 6500 23564 6502
rect 23620 6500 23644 6502
rect 23700 6500 23724 6502
rect 23780 6500 23786 6502
rect 23478 6480 23786 6500
rect 23478 5468 23786 5488
rect 23478 5466 23484 5468
rect 23540 5466 23564 5468
rect 23620 5466 23644 5468
rect 23700 5466 23724 5468
rect 23780 5466 23786 5468
rect 23540 5414 23542 5466
rect 23722 5414 23724 5466
rect 23478 5412 23484 5414
rect 23540 5412 23564 5414
rect 23620 5412 23644 5414
rect 23700 5412 23724 5414
rect 23780 5412 23786 5414
rect 23478 5392 23786 5412
rect 23478 4380 23786 4400
rect 23478 4378 23484 4380
rect 23540 4378 23564 4380
rect 23620 4378 23644 4380
rect 23700 4378 23724 4380
rect 23780 4378 23786 4380
rect 23540 4326 23542 4378
rect 23722 4326 23724 4378
rect 23478 4324 23484 4326
rect 23540 4324 23564 4326
rect 23620 4324 23644 4326
rect 23700 4324 23724 4326
rect 23780 4324 23786 4326
rect 23478 4304 23786 4324
rect 23478 3292 23786 3312
rect 23478 3290 23484 3292
rect 23540 3290 23564 3292
rect 23620 3290 23644 3292
rect 23700 3290 23724 3292
rect 23780 3290 23786 3292
rect 23540 3238 23542 3290
rect 23722 3238 23724 3290
rect 23478 3236 23484 3238
rect 23540 3236 23564 3238
rect 23620 3236 23644 3238
rect 23700 3236 23724 3238
rect 23780 3236 23786 3238
rect 23478 3216 23786 3236
rect 25148 3194 25176 25774
rect 25228 18148 25280 18154
rect 25228 18090 25280 18096
rect 22836 3188 22888 3194
rect 22836 3130 22888 3136
rect 25136 3188 25188 3194
rect 25136 3130 25188 3136
rect 22848 2446 22876 3130
rect 25148 3058 25176 3130
rect 25136 3052 25188 3058
rect 25136 2994 25188 3000
rect 24492 2848 24544 2854
rect 24492 2790 24544 2796
rect 22100 2440 22152 2446
rect 22100 2382 22152 2388
rect 22836 2440 22888 2446
rect 23480 2440 23532 2446
rect 22836 2382 22888 2388
rect 23216 2388 23480 2394
rect 23216 2382 23532 2388
rect 23216 2366 23520 2382
rect 22560 2304 22612 2310
rect 22560 2246 22612 2252
rect 22572 800 22600 2246
rect 23216 800 23244 2366
rect 23848 2304 23900 2310
rect 23848 2246 23900 2252
rect 23478 2204 23786 2224
rect 23478 2202 23484 2204
rect 23540 2202 23564 2204
rect 23620 2202 23644 2204
rect 23700 2202 23724 2204
rect 23780 2202 23786 2204
rect 23540 2150 23542 2202
rect 23722 2150 23724 2202
rect 23478 2148 23484 2150
rect 23540 2148 23564 2150
rect 23620 2148 23644 2150
rect 23700 2148 23724 2150
rect 23780 2148 23786 2150
rect 23478 2128 23786 2148
rect 23860 800 23888 2246
rect 24504 800 24532 2790
rect 25240 2446 25268 18090
rect 25504 17536 25556 17542
rect 25504 17478 25556 17484
rect 25516 3058 25544 17478
rect 25884 17338 25912 33458
rect 27264 33114 27292 35278
rect 28184 35278 28410 35306
rect 28184 33658 28212 35278
rect 28354 35200 28410 35278
rect 28998 35306 29054 36000
rect 29642 35306 29698 36000
rect 28998 35278 29132 35306
rect 28998 35200 29054 35278
rect 29104 33658 29132 35278
rect 29642 35278 29960 35306
rect 29642 35200 29698 35278
rect 29932 33658 29960 35278
rect 30286 35200 30342 36000
rect 30930 35306 30986 36000
rect 30760 35278 30986 35306
rect 28172 33652 28224 33658
rect 28172 33594 28224 33600
rect 29092 33652 29144 33658
rect 29092 33594 29144 33600
rect 29920 33652 29972 33658
rect 30300 33640 30328 35200
rect 30300 33612 30420 33640
rect 29920 33594 29972 33600
rect 30392 33522 30420 33612
rect 28724 33516 28776 33522
rect 28724 33458 28776 33464
rect 30380 33516 30432 33522
rect 30380 33458 30432 33464
rect 27344 33448 27396 33454
rect 27344 33390 27396 33396
rect 27620 33448 27672 33454
rect 27620 33390 27672 33396
rect 27252 33108 27304 33114
rect 27252 33050 27304 33056
rect 27252 18284 27304 18290
rect 27252 18226 27304 18232
rect 25872 17332 25924 17338
rect 25872 17274 25924 17280
rect 25504 3052 25556 3058
rect 25504 2994 25556 3000
rect 27068 2848 27120 2854
rect 27068 2790 27120 2796
rect 25228 2440 25280 2446
rect 25228 2382 25280 2388
rect 25136 2304 25188 2310
rect 25136 2246 25188 2252
rect 26424 2304 26476 2310
rect 26424 2246 26476 2252
rect 25148 800 25176 2246
rect 26436 800 26464 2246
rect 27080 800 27108 2790
rect 27264 2514 27292 18226
rect 27356 17678 27384 33390
rect 27632 18358 27660 33390
rect 27896 32904 27948 32910
rect 27896 32846 27948 32852
rect 27908 32502 27936 32846
rect 28736 32774 28764 33458
rect 29110 33212 29418 33232
rect 29110 33210 29116 33212
rect 29172 33210 29196 33212
rect 29252 33210 29276 33212
rect 29332 33210 29356 33212
rect 29412 33210 29418 33212
rect 29172 33158 29174 33210
rect 29354 33158 29356 33210
rect 29110 33156 29116 33158
rect 29172 33156 29196 33158
rect 29252 33156 29276 33158
rect 29332 33156 29356 33158
rect 29412 33156 29418 33158
rect 29110 33136 29418 33156
rect 30392 33114 30420 33458
rect 30760 33114 30788 35278
rect 30930 35200 30986 35278
rect 31574 35306 31630 36000
rect 32218 35306 32274 36000
rect 31574 35278 31708 35306
rect 31574 35200 31630 35278
rect 31680 33640 31708 35278
rect 32218 35278 32536 35306
rect 32218 35200 32274 35278
rect 31760 33652 31812 33658
rect 31680 33612 31760 33640
rect 31760 33594 31812 33600
rect 31208 33448 31260 33454
rect 31208 33390 31260 33396
rect 30840 33312 30892 33318
rect 30840 33254 30892 33260
rect 30380 33108 30432 33114
rect 30380 33050 30432 33056
rect 30748 33108 30800 33114
rect 30748 33050 30800 33056
rect 30760 32978 30788 33050
rect 29920 32972 29972 32978
rect 29920 32914 29972 32920
rect 30748 32972 30800 32978
rect 30748 32914 30800 32920
rect 28724 32768 28776 32774
rect 28724 32710 28776 32716
rect 28816 32768 28868 32774
rect 28816 32710 28868 32716
rect 27896 32496 27948 32502
rect 27896 32438 27948 32444
rect 28736 19242 28764 32710
rect 28828 32570 28856 32710
rect 28816 32564 28868 32570
rect 28816 32506 28868 32512
rect 29110 32124 29418 32144
rect 29110 32122 29116 32124
rect 29172 32122 29196 32124
rect 29252 32122 29276 32124
rect 29332 32122 29356 32124
rect 29412 32122 29418 32124
rect 29172 32070 29174 32122
rect 29354 32070 29356 32122
rect 29110 32068 29116 32070
rect 29172 32068 29196 32070
rect 29252 32068 29276 32070
rect 29332 32068 29356 32070
rect 29412 32068 29418 32070
rect 29110 32048 29418 32068
rect 29110 31036 29418 31056
rect 29110 31034 29116 31036
rect 29172 31034 29196 31036
rect 29252 31034 29276 31036
rect 29332 31034 29356 31036
rect 29412 31034 29418 31036
rect 29172 30982 29174 31034
rect 29354 30982 29356 31034
rect 29110 30980 29116 30982
rect 29172 30980 29196 30982
rect 29252 30980 29276 30982
rect 29332 30980 29356 30982
rect 29412 30980 29418 30982
rect 29110 30960 29418 30980
rect 29110 29948 29418 29968
rect 29110 29946 29116 29948
rect 29172 29946 29196 29948
rect 29252 29946 29276 29948
rect 29332 29946 29356 29948
rect 29412 29946 29418 29948
rect 29172 29894 29174 29946
rect 29354 29894 29356 29946
rect 29110 29892 29116 29894
rect 29172 29892 29196 29894
rect 29252 29892 29276 29894
rect 29332 29892 29356 29894
rect 29412 29892 29418 29894
rect 29110 29872 29418 29892
rect 29110 28860 29418 28880
rect 29110 28858 29116 28860
rect 29172 28858 29196 28860
rect 29252 28858 29276 28860
rect 29332 28858 29356 28860
rect 29412 28858 29418 28860
rect 29172 28806 29174 28858
rect 29354 28806 29356 28858
rect 29110 28804 29116 28806
rect 29172 28804 29196 28806
rect 29252 28804 29276 28806
rect 29332 28804 29356 28806
rect 29412 28804 29418 28806
rect 29110 28784 29418 28804
rect 29110 27772 29418 27792
rect 29110 27770 29116 27772
rect 29172 27770 29196 27772
rect 29252 27770 29276 27772
rect 29332 27770 29356 27772
rect 29412 27770 29418 27772
rect 29172 27718 29174 27770
rect 29354 27718 29356 27770
rect 29110 27716 29116 27718
rect 29172 27716 29196 27718
rect 29252 27716 29276 27718
rect 29332 27716 29356 27718
rect 29412 27716 29418 27718
rect 29110 27696 29418 27716
rect 29110 26684 29418 26704
rect 29110 26682 29116 26684
rect 29172 26682 29196 26684
rect 29252 26682 29276 26684
rect 29332 26682 29356 26684
rect 29412 26682 29418 26684
rect 29172 26630 29174 26682
rect 29354 26630 29356 26682
rect 29110 26628 29116 26630
rect 29172 26628 29196 26630
rect 29252 26628 29276 26630
rect 29332 26628 29356 26630
rect 29412 26628 29418 26630
rect 29110 26608 29418 26628
rect 29110 25596 29418 25616
rect 29110 25594 29116 25596
rect 29172 25594 29196 25596
rect 29252 25594 29276 25596
rect 29332 25594 29356 25596
rect 29412 25594 29418 25596
rect 29172 25542 29174 25594
rect 29354 25542 29356 25594
rect 29110 25540 29116 25542
rect 29172 25540 29196 25542
rect 29252 25540 29276 25542
rect 29332 25540 29356 25542
rect 29412 25540 29418 25542
rect 29110 25520 29418 25540
rect 29110 24508 29418 24528
rect 29110 24506 29116 24508
rect 29172 24506 29196 24508
rect 29252 24506 29276 24508
rect 29332 24506 29356 24508
rect 29412 24506 29418 24508
rect 29172 24454 29174 24506
rect 29354 24454 29356 24506
rect 29110 24452 29116 24454
rect 29172 24452 29196 24454
rect 29252 24452 29276 24454
rect 29332 24452 29356 24454
rect 29412 24452 29418 24454
rect 29110 24432 29418 24452
rect 29110 23420 29418 23440
rect 29110 23418 29116 23420
rect 29172 23418 29196 23420
rect 29252 23418 29276 23420
rect 29332 23418 29356 23420
rect 29412 23418 29418 23420
rect 29172 23366 29174 23418
rect 29354 23366 29356 23418
rect 29110 23364 29116 23366
rect 29172 23364 29196 23366
rect 29252 23364 29276 23366
rect 29332 23364 29356 23366
rect 29412 23364 29418 23366
rect 29110 23344 29418 23364
rect 29110 22332 29418 22352
rect 29110 22330 29116 22332
rect 29172 22330 29196 22332
rect 29252 22330 29276 22332
rect 29332 22330 29356 22332
rect 29412 22330 29418 22332
rect 29172 22278 29174 22330
rect 29354 22278 29356 22330
rect 29110 22276 29116 22278
rect 29172 22276 29196 22278
rect 29252 22276 29276 22278
rect 29332 22276 29356 22278
rect 29412 22276 29418 22278
rect 29110 22256 29418 22276
rect 29110 21244 29418 21264
rect 29110 21242 29116 21244
rect 29172 21242 29196 21244
rect 29252 21242 29276 21244
rect 29332 21242 29356 21244
rect 29412 21242 29418 21244
rect 29172 21190 29174 21242
rect 29354 21190 29356 21242
rect 29110 21188 29116 21190
rect 29172 21188 29196 21190
rect 29252 21188 29276 21190
rect 29332 21188 29356 21190
rect 29412 21188 29418 21190
rect 29110 21168 29418 21188
rect 29110 20156 29418 20176
rect 29110 20154 29116 20156
rect 29172 20154 29196 20156
rect 29252 20154 29276 20156
rect 29332 20154 29356 20156
rect 29412 20154 29418 20156
rect 29172 20102 29174 20154
rect 29354 20102 29356 20154
rect 29110 20100 29116 20102
rect 29172 20100 29196 20102
rect 29252 20100 29276 20102
rect 29332 20100 29356 20102
rect 29412 20100 29418 20102
rect 29110 20080 29418 20100
rect 28724 19236 28776 19242
rect 28724 19178 28776 19184
rect 29110 19068 29418 19088
rect 29110 19066 29116 19068
rect 29172 19066 29196 19068
rect 29252 19066 29276 19068
rect 29332 19066 29356 19068
rect 29412 19066 29418 19068
rect 29172 19014 29174 19066
rect 29354 19014 29356 19066
rect 29110 19012 29116 19014
rect 29172 19012 29196 19014
rect 29252 19012 29276 19014
rect 29332 19012 29356 19014
rect 29412 19012 29418 19014
rect 29110 18992 29418 19012
rect 29000 18828 29052 18834
rect 29000 18770 29052 18776
rect 29012 18426 29040 18770
rect 29184 18760 29236 18766
rect 29184 18702 29236 18708
rect 29196 18426 29224 18702
rect 29552 18624 29604 18630
rect 29552 18566 29604 18572
rect 29000 18420 29052 18426
rect 29000 18362 29052 18368
rect 29184 18420 29236 18426
rect 29184 18362 29236 18368
rect 29564 18358 29592 18566
rect 29932 18426 29960 32914
rect 30380 32428 30432 32434
rect 30380 32370 30432 32376
rect 30392 30802 30420 32370
rect 30380 30796 30432 30802
rect 30380 30738 30432 30744
rect 30852 28082 30880 33254
rect 30840 28076 30892 28082
rect 30840 28018 30892 28024
rect 29920 18420 29972 18426
rect 29920 18362 29972 18368
rect 30012 18420 30064 18426
rect 30012 18362 30064 18368
rect 27620 18352 27672 18358
rect 27620 18294 27672 18300
rect 29552 18352 29604 18358
rect 29552 18294 29604 18300
rect 29460 18284 29512 18290
rect 29460 18226 29512 18232
rect 29110 17980 29418 18000
rect 29110 17978 29116 17980
rect 29172 17978 29196 17980
rect 29252 17978 29276 17980
rect 29332 17978 29356 17980
rect 29412 17978 29418 17980
rect 29172 17926 29174 17978
rect 29354 17926 29356 17978
rect 29110 17924 29116 17926
rect 29172 17924 29196 17926
rect 29252 17924 29276 17926
rect 29332 17924 29356 17926
rect 29412 17924 29418 17926
rect 29110 17904 29418 17924
rect 27344 17672 27396 17678
rect 27344 17614 27396 17620
rect 29472 17202 29500 18226
rect 30024 18086 30052 18362
rect 31220 18358 31248 33390
rect 32312 33380 32364 33386
rect 32312 33322 32364 33328
rect 31944 32972 31996 32978
rect 31944 32914 31996 32920
rect 31300 32904 31352 32910
rect 31300 32846 31352 32852
rect 31312 26382 31340 32846
rect 31956 32230 31984 32914
rect 31944 32224 31996 32230
rect 31944 32166 31996 32172
rect 31300 26376 31352 26382
rect 31300 26318 31352 26324
rect 31852 25220 31904 25226
rect 31852 25162 31904 25168
rect 31864 22642 31892 25162
rect 31760 22636 31812 22642
rect 31760 22578 31812 22584
rect 31852 22636 31904 22642
rect 31852 22578 31904 22584
rect 31772 21554 31800 22578
rect 31760 21548 31812 21554
rect 31760 21490 31812 21496
rect 31760 19508 31812 19514
rect 31760 19450 31812 19456
rect 31772 18698 31800 19450
rect 31760 18692 31812 18698
rect 31760 18634 31812 18640
rect 31956 18426 31984 32166
rect 32324 26790 32352 33322
rect 32508 33114 32536 35278
rect 33506 35200 33562 36000
rect 33782 35456 33838 35465
rect 33612 35414 33782 35442
rect 33324 33516 33376 33522
rect 33324 33458 33376 33464
rect 33232 33448 33284 33454
rect 33138 33416 33194 33425
rect 32864 33380 32916 33386
rect 33232 33390 33284 33396
rect 33138 33351 33194 33360
rect 32864 33322 32916 33328
rect 32496 33108 32548 33114
rect 32496 33050 32548 33056
rect 32772 32836 32824 32842
rect 32772 32778 32824 32784
rect 32784 32570 32812 32778
rect 32772 32564 32824 32570
rect 32772 32506 32824 32512
rect 32312 26784 32364 26790
rect 32312 26726 32364 26732
rect 32496 26512 32548 26518
rect 32496 26454 32548 26460
rect 31944 18420 31996 18426
rect 31944 18362 31996 18368
rect 32508 18358 32536 26454
rect 31208 18352 31260 18358
rect 31208 18294 31260 18300
rect 32496 18352 32548 18358
rect 32496 18294 32548 18300
rect 32876 18290 32904 33322
rect 33152 33114 33180 33351
rect 33140 33108 33192 33114
rect 33140 33050 33192 33056
rect 32956 32904 33008 32910
rect 32956 32846 33008 32852
rect 32968 31822 32996 32846
rect 33244 32026 33272 33390
rect 33336 32366 33364 33458
rect 33520 32450 33548 35200
rect 33612 33454 33640 35414
rect 33782 35391 33838 35400
rect 34150 35200 34206 36000
rect 34794 35306 34850 36000
rect 34532 35278 34850 35306
rect 33690 34096 33746 34105
rect 33690 34031 33746 34040
rect 33600 33448 33652 33454
rect 33600 33390 33652 33396
rect 33704 33114 33732 34031
rect 33784 33448 33836 33454
rect 33784 33390 33836 33396
rect 33692 33108 33744 33114
rect 33692 33050 33744 33056
rect 33796 33046 33824 33390
rect 33784 33040 33836 33046
rect 33784 32982 33836 32988
rect 34164 32570 34192 35200
rect 34242 34776 34298 34785
rect 34242 34711 34298 34720
rect 34256 32910 34284 34711
rect 34428 33516 34480 33522
rect 34532 33504 34560 35278
rect 34794 35200 34850 35278
rect 35438 35200 35494 36000
rect 34480 33476 34560 33504
rect 34428 33458 34480 33464
rect 34244 32904 34296 32910
rect 34244 32846 34296 32852
rect 34152 32564 34204 32570
rect 34152 32506 34204 32512
rect 33428 32434 33548 32450
rect 33416 32428 33548 32434
rect 33468 32422 33548 32428
rect 33600 32428 33652 32434
rect 33416 32370 33468 32376
rect 33600 32370 33652 32376
rect 33324 32360 33376 32366
rect 33324 32302 33376 32308
rect 33428 32026 33456 32370
rect 33232 32020 33284 32026
rect 33232 31962 33284 31968
rect 33416 32020 33468 32026
rect 33416 31962 33468 31968
rect 33612 31906 33640 32370
rect 34244 32224 34296 32230
rect 34244 32166 34296 32172
rect 34256 32065 34284 32166
rect 34242 32056 34298 32065
rect 35452 32026 35480 35200
rect 34242 31991 34298 32000
rect 35440 32020 35492 32026
rect 35440 31962 35492 31968
rect 33428 31878 33640 31906
rect 32956 31816 33008 31822
rect 32956 31758 33008 31764
rect 30380 18284 30432 18290
rect 30380 18226 30432 18232
rect 32864 18284 32916 18290
rect 32864 18226 32916 18232
rect 30392 18086 30420 18226
rect 30932 18148 30984 18154
rect 30932 18090 30984 18096
rect 30012 18080 30064 18086
rect 30012 18022 30064 18028
rect 30380 18080 30432 18086
rect 30380 18022 30432 18028
rect 29460 17196 29512 17202
rect 29460 17138 29512 17144
rect 29828 17196 29880 17202
rect 29828 17138 29880 17144
rect 29110 16892 29418 16912
rect 29110 16890 29116 16892
rect 29172 16890 29196 16892
rect 29252 16890 29276 16892
rect 29332 16890 29356 16892
rect 29412 16890 29418 16892
rect 29172 16838 29174 16890
rect 29354 16838 29356 16890
rect 29110 16836 29116 16838
rect 29172 16836 29196 16838
rect 29252 16836 29276 16838
rect 29332 16836 29356 16838
rect 29412 16836 29418 16838
rect 29110 16816 29418 16836
rect 29110 15804 29418 15824
rect 29110 15802 29116 15804
rect 29172 15802 29196 15804
rect 29252 15802 29276 15804
rect 29332 15802 29356 15804
rect 29412 15802 29418 15804
rect 29172 15750 29174 15802
rect 29354 15750 29356 15802
rect 29110 15748 29116 15750
rect 29172 15748 29196 15750
rect 29252 15748 29276 15750
rect 29332 15748 29356 15750
rect 29412 15748 29418 15750
rect 29110 15728 29418 15748
rect 29110 14716 29418 14736
rect 29110 14714 29116 14716
rect 29172 14714 29196 14716
rect 29252 14714 29276 14716
rect 29332 14714 29356 14716
rect 29412 14714 29418 14716
rect 29172 14662 29174 14714
rect 29354 14662 29356 14714
rect 29110 14660 29116 14662
rect 29172 14660 29196 14662
rect 29252 14660 29276 14662
rect 29332 14660 29356 14662
rect 29412 14660 29418 14662
rect 29110 14640 29418 14660
rect 29110 13628 29418 13648
rect 29110 13626 29116 13628
rect 29172 13626 29196 13628
rect 29252 13626 29276 13628
rect 29332 13626 29356 13628
rect 29412 13626 29418 13628
rect 29172 13574 29174 13626
rect 29354 13574 29356 13626
rect 29110 13572 29116 13574
rect 29172 13572 29196 13574
rect 29252 13572 29276 13574
rect 29332 13572 29356 13574
rect 29412 13572 29418 13574
rect 29110 13552 29418 13572
rect 29110 12540 29418 12560
rect 29110 12538 29116 12540
rect 29172 12538 29196 12540
rect 29252 12538 29276 12540
rect 29332 12538 29356 12540
rect 29412 12538 29418 12540
rect 29172 12486 29174 12538
rect 29354 12486 29356 12538
rect 29110 12484 29116 12486
rect 29172 12484 29196 12486
rect 29252 12484 29276 12486
rect 29332 12484 29356 12486
rect 29412 12484 29418 12486
rect 29110 12464 29418 12484
rect 29110 11452 29418 11472
rect 29110 11450 29116 11452
rect 29172 11450 29196 11452
rect 29252 11450 29276 11452
rect 29332 11450 29356 11452
rect 29412 11450 29418 11452
rect 29172 11398 29174 11450
rect 29354 11398 29356 11450
rect 29110 11396 29116 11398
rect 29172 11396 29196 11398
rect 29252 11396 29276 11398
rect 29332 11396 29356 11398
rect 29412 11396 29418 11398
rect 29110 11376 29418 11396
rect 29110 10364 29418 10384
rect 29110 10362 29116 10364
rect 29172 10362 29196 10364
rect 29252 10362 29276 10364
rect 29332 10362 29356 10364
rect 29412 10362 29418 10364
rect 29172 10310 29174 10362
rect 29354 10310 29356 10362
rect 29110 10308 29116 10310
rect 29172 10308 29196 10310
rect 29252 10308 29276 10310
rect 29332 10308 29356 10310
rect 29412 10308 29418 10310
rect 29110 10288 29418 10308
rect 29110 9276 29418 9296
rect 29110 9274 29116 9276
rect 29172 9274 29196 9276
rect 29252 9274 29276 9276
rect 29332 9274 29356 9276
rect 29412 9274 29418 9276
rect 29172 9222 29174 9274
rect 29354 9222 29356 9274
rect 29110 9220 29116 9222
rect 29172 9220 29196 9222
rect 29252 9220 29276 9222
rect 29332 9220 29356 9222
rect 29412 9220 29418 9222
rect 29110 9200 29418 9220
rect 29110 8188 29418 8208
rect 29110 8186 29116 8188
rect 29172 8186 29196 8188
rect 29252 8186 29276 8188
rect 29332 8186 29356 8188
rect 29412 8186 29418 8188
rect 29172 8134 29174 8186
rect 29354 8134 29356 8186
rect 29110 8132 29116 8134
rect 29172 8132 29196 8134
rect 29252 8132 29276 8134
rect 29332 8132 29356 8134
rect 29412 8132 29418 8134
rect 29110 8112 29418 8132
rect 29110 7100 29418 7120
rect 29110 7098 29116 7100
rect 29172 7098 29196 7100
rect 29252 7098 29276 7100
rect 29332 7098 29356 7100
rect 29412 7098 29418 7100
rect 29172 7046 29174 7098
rect 29354 7046 29356 7098
rect 29110 7044 29116 7046
rect 29172 7044 29196 7046
rect 29252 7044 29276 7046
rect 29332 7044 29356 7046
rect 29412 7044 29418 7046
rect 29110 7024 29418 7044
rect 29110 6012 29418 6032
rect 29110 6010 29116 6012
rect 29172 6010 29196 6012
rect 29252 6010 29276 6012
rect 29332 6010 29356 6012
rect 29412 6010 29418 6012
rect 29172 5958 29174 6010
rect 29354 5958 29356 6010
rect 29110 5956 29116 5958
rect 29172 5956 29196 5958
rect 29252 5956 29276 5958
rect 29332 5956 29356 5958
rect 29412 5956 29418 5958
rect 29110 5936 29418 5956
rect 29110 4924 29418 4944
rect 29110 4922 29116 4924
rect 29172 4922 29196 4924
rect 29252 4922 29276 4924
rect 29332 4922 29356 4924
rect 29412 4922 29418 4924
rect 29172 4870 29174 4922
rect 29354 4870 29356 4922
rect 29110 4868 29116 4870
rect 29172 4868 29196 4870
rect 29252 4868 29276 4870
rect 29332 4868 29356 4870
rect 29412 4868 29418 4870
rect 29110 4848 29418 4868
rect 29110 3836 29418 3856
rect 29110 3834 29116 3836
rect 29172 3834 29196 3836
rect 29252 3834 29276 3836
rect 29332 3834 29356 3836
rect 29412 3834 29418 3836
rect 29172 3782 29174 3834
rect 29354 3782 29356 3834
rect 29110 3780 29116 3782
rect 29172 3780 29196 3782
rect 29252 3780 29276 3782
rect 29332 3780 29356 3782
rect 29412 3780 29418 3782
rect 29110 3760 29418 3780
rect 29736 3528 29788 3534
rect 29736 3470 29788 3476
rect 29748 3194 29776 3470
rect 29736 3188 29788 3194
rect 29736 3130 29788 3136
rect 28632 3120 28684 3126
rect 28632 3062 28684 3068
rect 28080 2984 28132 2990
rect 28080 2926 28132 2932
rect 27252 2508 27304 2514
rect 27252 2450 27304 2456
rect 28092 2446 28120 2926
rect 28644 2650 28672 3062
rect 29644 3052 29696 3058
rect 29644 2994 29696 3000
rect 29460 2848 29512 2854
rect 29460 2790 29512 2796
rect 29110 2748 29418 2768
rect 29110 2746 29116 2748
rect 29172 2746 29196 2748
rect 29252 2746 29276 2748
rect 29332 2746 29356 2748
rect 29412 2746 29418 2748
rect 29172 2694 29174 2746
rect 29354 2694 29356 2746
rect 29110 2692 29116 2694
rect 29172 2692 29196 2694
rect 29252 2692 29276 2694
rect 29332 2692 29356 2694
rect 29412 2692 29418 2694
rect 29110 2672 29418 2692
rect 28632 2644 28684 2650
rect 28632 2586 28684 2592
rect 29472 2446 29500 2790
rect 28080 2440 28132 2446
rect 28080 2382 28132 2388
rect 28356 2440 28408 2446
rect 28356 2382 28408 2388
rect 29000 2440 29052 2446
rect 29000 2382 29052 2388
rect 29460 2440 29512 2446
rect 29460 2382 29512 2388
rect 27712 2304 27764 2310
rect 27712 2246 27764 2252
rect 27724 800 27752 2246
rect 28368 800 28396 2382
rect 29012 800 29040 2382
rect 29656 800 29684 2994
rect 29840 2514 29868 17138
rect 30104 5160 30156 5166
rect 30104 5102 30156 5108
rect 30116 4690 30144 5102
rect 30104 4684 30156 4690
rect 30104 4626 30156 4632
rect 30392 3126 30420 18022
rect 30380 3120 30432 3126
rect 30380 3062 30432 3068
rect 29828 2508 29880 2514
rect 29828 2450 29880 2456
rect 30944 2446 30972 18090
rect 31300 18080 31352 18086
rect 31300 18022 31352 18028
rect 31312 3058 31340 18022
rect 32968 17898 32996 31758
rect 33428 31142 33456 31878
rect 33600 31816 33652 31822
rect 33600 31758 33652 31764
rect 33416 31136 33468 31142
rect 33416 31078 33468 31084
rect 33048 25424 33100 25430
rect 33048 25366 33100 25372
rect 33060 23322 33088 25366
rect 33048 23316 33100 23322
rect 33048 23258 33100 23264
rect 33428 18834 33456 31078
rect 33612 29850 33640 31758
rect 34334 31376 34390 31385
rect 34334 31311 34336 31320
rect 34388 31311 34390 31320
rect 34336 31282 34388 31288
rect 33692 31136 33744 31142
rect 33692 31078 33744 31084
rect 33600 29844 33652 29850
rect 33600 29786 33652 29792
rect 33508 20936 33560 20942
rect 33508 20878 33560 20884
rect 33520 20505 33548 20878
rect 33506 20496 33562 20505
rect 33506 20431 33562 20440
rect 33416 18828 33468 18834
rect 33416 18770 33468 18776
rect 33704 18290 33732 31078
rect 34060 30932 34112 30938
rect 34060 30874 34112 30880
rect 33876 30048 33928 30054
rect 33876 29990 33928 29996
rect 33888 29170 33916 29990
rect 34072 29170 34100 30874
rect 34336 30728 34388 30734
rect 34334 30696 34336 30705
rect 34388 30696 34390 30705
rect 34334 30631 34390 30640
rect 34348 30394 34376 30631
rect 34336 30388 34388 30394
rect 34336 30330 34388 30336
rect 34336 30252 34388 30258
rect 34336 30194 34388 30200
rect 34348 30025 34376 30194
rect 34334 30016 34390 30025
rect 34334 29951 34390 29960
rect 34336 29640 34388 29646
rect 34336 29582 34388 29588
rect 34348 29345 34376 29582
rect 34334 29336 34390 29345
rect 34334 29271 34390 29280
rect 33876 29164 33928 29170
rect 33876 29106 33928 29112
rect 34060 29164 34112 29170
rect 34060 29106 34112 29112
rect 34072 29050 34100 29106
rect 33980 29022 34100 29050
rect 34244 29028 34296 29034
rect 33980 28762 34008 29022
rect 34244 28970 34296 28976
rect 34060 28960 34112 28966
rect 34060 28902 34112 28908
rect 33968 28756 34020 28762
rect 33968 28698 34020 28704
rect 34072 28082 34100 28902
rect 34256 28665 34284 28970
rect 34242 28656 34298 28665
rect 34242 28591 34298 28600
rect 34060 28076 34112 28082
rect 34060 28018 34112 28024
rect 34242 27976 34298 27985
rect 34242 27911 34244 27920
rect 34296 27911 34298 27920
rect 34244 27882 34296 27888
rect 34060 27872 34112 27878
rect 34060 27814 34112 27820
rect 34072 25294 34100 27814
rect 34244 26988 34296 26994
rect 34244 26930 34296 26936
rect 34152 26784 34204 26790
rect 34152 26726 34204 26732
rect 34060 25288 34112 25294
rect 34060 25230 34112 25236
rect 34060 24812 34112 24818
rect 34060 24754 34112 24760
rect 33876 24132 33928 24138
rect 33876 24074 33928 24080
rect 33692 18284 33744 18290
rect 33692 18226 33744 18232
rect 32876 17870 32996 17898
rect 32876 17746 32904 17870
rect 32956 17808 33008 17814
rect 32956 17750 33008 17756
rect 32864 17740 32916 17746
rect 32864 17682 32916 17688
rect 32404 17604 32456 17610
rect 32404 17546 32456 17552
rect 31760 16040 31812 16046
rect 31760 15982 31812 15988
rect 31772 15094 31800 15982
rect 31760 15088 31812 15094
rect 31760 15030 31812 15036
rect 32416 7410 32444 17546
rect 32404 7404 32456 7410
rect 32404 7346 32456 7352
rect 31852 3528 31904 3534
rect 32404 3528 32456 3534
rect 31852 3470 31904 3476
rect 32402 3496 32404 3505
rect 32456 3496 32458 3505
rect 31300 3052 31352 3058
rect 31300 2994 31352 3000
rect 31864 2514 31892 3470
rect 32402 3431 32458 3440
rect 32416 3058 32444 3431
rect 32404 3052 32456 3058
rect 32404 2994 32456 3000
rect 32404 2916 32456 2922
rect 32404 2858 32456 2864
rect 32220 2848 32272 2854
rect 32220 2790 32272 2796
rect 31852 2508 31904 2514
rect 31852 2450 31904 2456
rect 30932 2440 30984 2446
rect 30932 2382 30984 2388
rect 31576 2440 31628 2446
rect 31576 2382 31628 2388
rect 30288 2304 30340 2310
rect 30288 2246 30340 2252
rect 30300 800 30328 2246
rect 31588 800 31616 2382
rect 32232 800 32260 2790
rect 32416 2446 32444 2858
rect 32864 2848 32916 2854
rect 32864 2790 32916 2796
rect 32404 2440 32456 2446
rect 32404 2382 32456 2388
rect 32588 2304 32640 2310
rect 32588 2246 32640 2252
rect 32600 2145 32628 2246
rect 32586 2136 32642 2145
rect 32586 2071 32642 2080
rect 32876 800 32904 2790
rect 32968 2582 32996 17750
rect 33600 17196 33652 17202
rect 33600 17138 33652 17144
rect 33140 17128 33192 17134
rect 33140 17070 33192 17076
rect 33152 13938 33180 17070
rect 33140 13932 33192 13938
rect 33140 13874 33192 13880
rect 33612 10266 33640 17138
rect 33692 13184 33744 13190
rect 33692 13126 33744 13132
rect 33600 10260 33652 10266
rect 33600 10202 33652 10208
rect 33704 9926 33732 13126
rect 33692 9920 33744 9926
rect 33692 9862 33744 9868
rect 33888 4146 33916 24074
rect 34072 20602 34100 24754
rect 34164 24138 34192 26726
rect 34256 26625 34284 26930
rect 34242 26616 34298 26625
rect 34242 26551 34298 26560
rect 34336 26376 34388 26382
rect 34336 26318 34388 26324
rect 34348 25945 34376 26318
rect 34334 25936 34390 25945
rect 34334 25871 34390 25880
rect 34242 25256 34298 25265
rect 34242 25191 34298 25200
rect 34256 25158 34284 25191
rect 34244 25152 34296 25158
rect 34244 25094 34296 25100
rect 34244 24608 34296 24614
rect 34242 24576 34244 24585
rect 34296 24576 34298 24585
rect 34242 24511 34298 24520
rect 34152 24132 34204 24138
rect 34152 24074 34204 24080
rect 34242 23896 34298 23905
rect 34242 23831 34298 23840
rect 34256 23798 34284 23831
rect 34244 23792 34296 23798
rect 34244 23734 34296 23740
rect 34244 23248 34296 23254
rect 34242 23216 34244 23225
rect 34296 23216 34298 23225
rect 34242 23151 34298 23160
rect 34336 22568 34388 22574
rect 34334 22536 34336 22545
rect 34388 22536 34390 22545
rect 34334 22471 34390 22480
rect 34348 22234 34376 22471
rect 34336 22228 34388 22234
rect 34336 22170 34388 22176
rect 34336 21888 34388 21894
rect 34336 21830 34388 21836
rect 34348 21486 34376 21830
rect 34336 21480 34388 21486
rect 34336 21422 34388 21428
rect 34348 21185 34376 21422
rect 34334 21176 34390 21185
rect 34334 21111 34390 21120
rect 34060 20596 34112 20602
rect 34060 20538 34112 20544
rect 34152 20460 34204 20466
rect 34152 20402 34204 20408
rect 34164 20058 34192 20402
rect 34152 20052 34204 20058
rect 34152 19994 34204 20000
rect 34336 19848 34388 19854
rect 34334 19816 34336 19825
rect 34388 19816 34390 19825
rect 34334 19751 34390 19760
rect 34336 19372 34388 19378
rect 34336 19314 34388 19320
rect 34348 19145 34376 19314
rect 34334 19136 34390 19145
rect 34334 19071 34390 19080
rect 34336 18760 34388 18766
rect 34336 18702 34388 18708
rect 34348 18465 34376 18702
rect 34334 18456 34390 18465
rect 34334 18391 34390 18400
rect 34060 18284 34112 18290
rect 34060 18226 34112 18232
rect 33968 18080 34020 18086
rect 33968 18022 34020 18028
rect 33980 7886 34008 18022
rect 34072 17338 34100 18226
rect 34244 18080 34296 18086
rect 34244 18022 34296 18028
rect 34256 17785 34284 18022
rect 34242 17776 34298 17785
rect 34242 17711 34298 17720
rect 34060 17332 34112 17338
rect 34060 17274 34112 17280
rect 34242 17096 34298 17105
rect 34242 17031 34244 17040
rect 34296 17031 34298 17040
rect 34244 17002 34296 17008
rect 34336 16448 34388 16454
rect 34336 16390 34388 16396
rect 34348 16046 34376 16390
rect 34336 16040 34388 16046
rect 34336 15982 34388 15988
rect 34348 15745 34376 15982
rect 34334 15736 34390 15745
rect 34334 15671 34390 15680
rect 34060 15496 34112 15502
rect 34060 15438 34112 15444
rect 34072 15162 34100 15438
rect 34244 15360 34296 15366
rect 34244 15302 34296 15308
rect 34060 15156 34112 15162
rect 34060 15098 34112 15104
rect 34256 15065 34284 15302
rect 34242 15056 34298 15065
rect 34152 15020 34204 15026
rect 34242 14991 34298 15000
rect 34152 14962 34204 14968
rect 34164 14618 34192 14962
rect 34152 14612 34204 14618
rect 34152 14554 34204 14560
rect 34336 14408 34388 14414
rect 34334 14376 34336 14385
rect 34388 14376 34390 14385
rect 34334 14311 34390 14320
rect 34336 14272 34388 14278
rect 34336 14214 34388 14220
rect 34348 13870 34376 14214
rect 34336 13864 34388 13870
rect 34336 13806 34388 13812
rect 34348 13705 34376 13806
rect 34334 13696 34390 13705
rect 34334 13631 34390 13640
rect 34244 13184 34296 13190
rect 34244 13126 34296 13132
rect 34256 13025 34284 13126
rect 34242 13016 34298 13025
rect 34242 12951 34298 12960
rect 34244 12640 34296 12646
rect 34244 12582 34296 12588
rect 34256 12345 34284 12582
rect 34242 12336 34298 12345
rect 34242 12271 34298 12280
rect 34242 11656 34298 11665
rect 34242 11591 34244 11600
rect 34296 11591 34298 11600
rect 34244 11562 34296 11568
rect 34336 10056 34388 10062
rect 34336 9998 34388 10004
rect 34348 9625 34376 9998
rect 34334 9616 34390 9625
rect 34334 9551 34390 9560
rect 34242 8936 34298 8945
rect 34242 8871 34298 8880
rect 34256 8838 34284 8871
rect 34244 8832 34296 8838
rect 34244 8774 34296 8780
rect 34244 8492 34296 8498
rect 34244 8434 34296 8440
rect 34256 8265 34284 8434
rect 34242 8256 34298 8265
rect 34242 8191 34298 8200
rect 33968 7880 34020 7886
rect 33968 7822 34020 7828
rect 34244 7744 34296 7750
rect 34244 7686 34296 7692
rect 34256 7585 34284 7686
rect 34242 7576 34298 7585
rect 34242 7511 34298 7520
rect 34244 7200 34296 7206
rect 34244 7142 34296 7148
rect 34256 6905 34284 7142
rect 34242 6896 34298 6905
rect 34242 6831 34298 6840
rect 34244 6316 34296 6322
rect 34244 6258 34296 6264
rect 34256 6225 34284 6258
rect 34242 6216 34298 6225
rect 34242 6151 34298 6160
rect 34336 5568 34388 5574
rect 34336 5510 34388 5516
rect 34348 5166 34376 5510
rect 34336 5160 34388 5166
rect 34336 5102 34388 5108
rect 34348 4865 34376 5102
rect 34334 4856 34390 4865
rect 34334 4791 34390 4800
rect 34244 4480 34296 4486
rect 34244 4422 34296 4428
rect 34256 4185 34284 4422
rect 34242 4176 34298 4185
rect 33876 4140 33928 4146
rect 34242 4111 34298 4120
rect 33876 4082 33928 4088
rect 33876 3936 33928 3942
rect 33876 3878 33928 3884
rect 34244 3936 34296 3942
rect 34244 3878 34296 3884
rect 33140 3392 33192 3398
rect 33140 3334 33192 3340
rect 32956 2576 33008 2582
rect 32956 2518 33008 2524
rect 33152 2378 33180 3334
rect 33508 2984 33560 2990
rect 33508 2926 33560 2932
rect 33140 2372 33192 2378
rect 33140 2314 33192 2320
rect 33152 1465 33180 2314
rect 33138 1456 33194 1465
rect 33138 1391 33194 1400
rect 33520 800 33548 2926
rect 33888 2514 33916 3878
rect 34256 2825 34284 3878
rect 34520 3732 34572 3738
rect 34520 3674 34572 3680
rect 34532 3466 34560 3674
rect 34796 3664 34848 3670
rect 34796 3606 34848 3612
rect 34520 3460 34572 3466
rect 34520 3402 34572 3408
rect 34242 2816 34298 2825
rect 34242 2751 34298 2760
rect 33876 2508 33928 2514
rect 33876 2450 33928 2456
rect 3018 734 3096 762
rect 2962 711 3018 720
rect 3238 0 3294 800
rect 3882 0 3938 800
rect 4526 0 4582 800
rect 5814 0 5870 800
rect 6458 0 6514 800
rect 7102 0 7158 800
rect 7746 0 7802 800
rect 8390 0 8446 800
rect 9034 0 9090 800
rect 9678 0 9734 800
rect 10966 0 11022 800
rect 11610 0 11666 800
rect 12254 0 12310 800
rect 12898 0 12954 800
rect 13542 0 13598 800
rect 14186 0 14242 800
rect 14830 0 14886 800
rect 16118 0 16174 800
rect 16762 0 16818 800
rect 17406 0 17462 800
rect 18050 0 18106 800
rect 18694 0 18750 800
rect 19338 0 19394 800
rect 19982 0 20038 800
rect 21270 0 21326 800
rect 21914 0 21970 800
rect 22558 0 22614 800
rect 23202 0 23258 800
rect 23846 0 23902 800
rect 24490 0 24546 800
rect 25134 0 25190 800
rect 26422 0 26478 800
rect 27066 0 27122 800
rect 27710 0 27766 800
rect 28354 0 28410 800
rect 28998 0 29054 800
rect 29642 0 29698 800
rect 30286 0 30342 800
rect 31574 0 31630 800
rect 32218 0 32274 800
rect 32862 0 32918 800
rect 33506 0 33562 800
rect 33888 785 33916 2450
rect 34808 800 34836 3606
rect 35440 3460 35492 3466
rect 35440 3402 35492 3408
rect 35452 800 35480 3402
rect 33874 776 33930 785
rect 33874 711 33930 720
rect 34150 0 34206 800
rect 34794 0 34850 800
rect 35438 0 35494 800
<< via2 >>
rect 2962 35400 3018 35456
rect 2134 34040 2190 34096
rect 2870 34720 2926 34776
rect 1398 32000 1454 32056
rect 1674 31864 1730 31920
rect 1490 31320 1546 31376
rect 1490 30640 1546 30696
rect 1490 29280 1546 29336
rect 1674 28600 1730 28656
rect 1490 27940 1546 27976
rect 1490 27920 1492 27940
rect 1492 27920 1544 27940
rect 1544 27920 1546 27940
rect 1398 25880 1454 25936
rect 1490 24556 1492 24576
rect 1492 24556 1544 24576
rect 1544 24556 1546 24576
rect 1490 24520 1546 24556
rect 1490 23840 1546 23896
rect 1490 23160 1546 23216
rect 1490 22500 1546 22536
rect 1490 22480 1492 22500
rect 1492 22480 1544 22500
rect 1544 22480 1546 22500
rect 1490 21120 1546 21176
rect 1398 19796 1400 19816
rect 1400 19796 1452 19816
rect 1452 19796 1454 19816
rect 1398 19760 1454 19796
rect 1398 19080 1454 19136
rect 1490 17720 1546 17776
rect 1490 17060 1546 17096
rect 1490 17040 1492 17060
rect 1492 17040 1544 17060
rect 1544 17040 1546 17060
rect 1490 15680 1546 15736
rect 1398 15000 1454 15056
rect 1490 14320 1546 14376
rect 1490 12280 1546 12336
rect 1398 11636 1400 11656
rect 1400 11636 1452 11656
rect 1452 11636 1454 11656
rect 1398 11600 1454 11636
rect 1950 29960 2006 30016
rect 1674 12960 1730 13016
rect 1398 10240 1454 10296
rect 1490 8880 1546 8936
rect 1490 7520 1546 7576
rect 1490 6840 1546 6896
rect 1490 6180 1546 6216
rect 1490 6160 1492 6180
rect 1492 6160 1544 6180
rect 1544 6160 1546 6180
rect 1490 4800 1546 4856
rect 2134 18400 2190 18456
rect 6588 33210 6644 33212
rect 6668 33210 6724 33212
rect 6748 33210 6804 33212
rect 6828 33210 6884 33212
rect 6588 33158 6634 33210
rect 6634 33158 6644 33210
rect 6668 33158 6698 33210
rect 6698 33158 6710 33210
rect 6710 33158 6724 33210
rect 6748 33158 6762 33210
rect 6762 33158 6774 33210
rect 6774 33158 6804 33210
rect 6828 33158 6838 33210
rect 6838 33158 6884 33210
rect 6588 33156 6644 33158
rect 6668 33156 6724 33158
rect 6748 33156 6804 33158
rect 6828 33156 6884 33158
rect 6588 32122 6644 32124
rect 6668 32122 6724 32124
rect 6748 32122 6804 32124
rect 6828 32122 6884 32124
rect 6588 32070 6634 32122
rect 6634 32070 6644 32122
rect 6668 32070 6698 32122
rect 6698 32070 6710 32122
rect 6710 32070 6724 32122
rect 6748 32070 6762 32122
rect 6762 32070 6774 32122
rect 6774 32070 6804 32122
rect 6828 32070 6838 32122
rect 6838 32070 6884 32122
rect 6588 32068 6644 32070
rect 6668 32068 6724 32070
rect 6748 32068 6804 32070
rect 6828 32068 6884 32070
rect 6588 31034 6644 31036
rect 6668 31034 6724 31036
rect 6748 31034 6804 31036
rect 6828 31034 6884 31036
rect 6588 30982 6634 31034
rect 6634 30982 6644 31034
rect 6668 30982 6698 31034
rect 6698 30982 6710 31034
rect 6710 30982 6724 31034
rect 6748 30982 6762 31034
rect 6762 30982 6774 31034
rect 6774 30982 6804 31034
rect 6828 30982 6838 31034
rect 6838 30982 6884 31034
rect 6588 30980 6644 30982
rect 6668 30980 6724 30982
rect 6748 30980 6804 30982
rect 6828 30980 6884 30982
rect 6588 29946 6644 29948
rect 6668 29946 6724 29948
rect 6748 29946 6804 29948
rect 6828 29946 6884 29948
rect 6588 29894 6634 29946
rect 6634 29894 6644 29946
rect 6668 29894 6698 29946
rect 6698 29894 6710 29946
rect 6710 29894 6724 29946
rect 6748 29894 6762 29946
rect 6762 29894 6774 29946
rect 6774 29894 6804 29946
rect 6828 29894 6838 29946
rect 6838 29894 6884 29946
rect 6588 29892 6644 29894
rect 6668 29892 6724 29894
rect 6748 29892 6804 29894
rect 6828 29892 6884 29894
rect 6588 28858 6644 28860
rect 6668 28858 6724 28860
rect 6748 28858 6804 28860
rect 6828 28858 6884 28860
rect 6588 28806 6634 28858
rect 6634 28806 6644 28858
rect 6668 28806 6698 28858
rect 6698 28806 6710 28858
rect 6710 28806 6724 28858
rect 6748 28806 6762 28858
rect 6762 28806 6774 28858
rect 6774 28806 6804 28858
rect 6828 28806 6838 28858
rect 6838 28806 6884 28858
rect 6588 28804 6644 28806
rect 6668 28804 6724 28806
rect 6748 28804 6804 28806
rect 6828 28804 6884 28806
rect 6588 27770 6644 27772
rect 6668 27770 6724 27772
rect 6748 27770 6804 27772
rect 6828 27770 6884 27772
rect 6588 27718 6634 27770
rect 6634 27718 6644 27770
rect 6668 27718 6698 27770
rect 6698 27718 6710 27770
rect 6710 27718 6724 27770
rect 6748 27718 6762 27770
rect 6762 27718 6774 27770
rect 6774 27718 6804 27770
rect 6828 27718 6838 27770
rect 6838 27718 6884 27770
rect 6588 27716 6644 27718
rect 6668 27716 6724 27718
rect 6748 27716 6804 27718
rect 6828 27716 6884 27718
rect 6588 26682 6644 26684
rect 6668 26682 6724 26684
rect 6748 26682 6804 26684
rect 6828 26682 6884 26684
rect 6588 26630 6634 26682
rect 6634 26630 6644 26682
rect 6668 26630 6698 26682
rect 6698 26630 6710 26682
rect 6710 26630 6724 26682
rect 6748 26630 6762 26682
rect 6762 26630 6774 26682
rect 6774 26630 6804 26682
rect 6828 26630 6838 26682
rect 6838 26630 6884 26682
rect 6588 26628 6644 26630
rect 6668 26628 6724 26630
rect 6748 26628 6804 26630
rect 6828 26628 6884 26630
rect 6588 25594 6644 25596
rect 6668 25594 6724 25596
rect 6748 25594 6804 25596
rect 6828 25594 6884 25596
rect 6588 25542 6634 25594
rect 6634 25542 6644 25594
rect 6668 25542 6698 25594
rect 6698 25542 6710 25594
rect 6710 25542 6724 25594
rect 6748 25542 6762 25594
rect 6762 25542 6774 25594
rect 6774 25542 6804 25594
rect 6828 25542 6838 25594
rect 6838 25542 6884 25594
rect 6588 25540 6644 25542
rect 6668 25540 6724 25542
rect 6748 25540 6804 25542
rect 6828 25540 6884 25542
rect 6588 24506 6644 24508
rect 6668 24506 6724 24508
rect 6748 24506 6804 24508
rect 6828 24506 6884 24508
rect 6588 24454 6634 24506
rect 6634 24454 6644 24506
rect 6668 24454 6698 24506
rect 6698 24454 6710 24506
rect 6710 24454 6724 24506
rect 6748 24454 6762 24506
rect 6762 24454 6774 24506
rect 6774 24454 6804 24506
rect 6828 24454 6838 24506
rect 6838 24454 6884 24506
rect 6588 24452 6644 24454
rect 6668 24452 6724 24454
rect 6748 24452 6804 24454
rect 6828 24452 6884 24454
rect 6588 23418 6644 23420
rect 6668 23418 6724 23420
rect 6748 23418 6804 23420
rect 6828 23418 6884 23420
rect 6588 23366 6634 23418
rect 6634 23366 6644 23418
rect 6668 23366 6698 23418
rect 6698 23366 6710 23418
rect 6710 23366 6724 23418
rect 6748 23366 6762 23418
rect 6762 23366 6774 23418
rect 6774 23366 6804 23418
rect 6828 23366 6838 23418
rect 6838 23366 6884 23418
rect 6588 23364 6644 23366
rect 6668 23364 6724 23366
rect 6748 23364 6804 23366
rect 6828 23364 6884 23366
rect 6588 22330 6644 22332
rect 6668 22330 6724 22332
rect 6748 22330 6804 22332
rect 6828 22330 6884 22332
rect 6588 22278 6634 22330
rect 6634 22278 6644 22330
rect 6668 22278 6698 22330
rect 6698 22278 6710 22330
rect 6710 22278 6724 22330
rect 6748 22278 6762 22330
rect 6762 22278 6774 22330
rect 6774 22278 6804 22330
rect 6828 22278 6838 22330
rect 6838 22278 6884 22330
rect 6588 22276 6644 22278
rect 6668 22276 6724 22278
rect 6748 22276 6804 22278
rect 6828 22276 6884 22278
rect 6588 21242 6644 21244
rect 6668 21242 6724 21244
rect 6748 21242 6804 21244
rect 6828 21242 6884 21244
rect 6588 21190 6634 21242
rect 6634 21190 6644 21242
rect 6668 21190 6698 21242
rect 6698 21190 6710 21242
rect 6710 21190 6724 21242
rect 6748 21190 6762 21242
rect 6762 21190 6774 21242
rect 6774 21190 6804 21242
rect 6828 21190 6838 21242
rect 6838 21190 6884 21242
rect 6588 21188 6644 21190
rect 6668 21188 6724 21190
rect 6748 21188 6804 21190
rect 6828 21188 6884 21190
rect 6588 20154 6644 20156
rect 6668 20154 6724 20156
rect 6748 20154 6804 20156
rect 6828 20154 6884 20156
rect 6588 20102 6634 20154
rect 6634 20102 6644 20154
rect 6668 20102 6698 20154
rect 6698 20102 6710 20154
rect 6710 20102 6724 20154
rect 6748 20102 6762 20154
rect 6762 20102 6774 20154
rect 6774 20102 6804 20154
rect 6828 20102 6838 20154
rect 6838 20102 6884 20154
rect 6588 20100 6644 20102
rect 6668 20100 6724 20102
rect 6748 20100 6804 20102
rect 6828 20100 6884 20102
rect 6588 19066 6644 19068
rect 6668 19066 6724 19068
rect 6748 19066 6804 19068
rect 6828 19066 6884 19068
rect 6588 19014 6634 19066
rect 6634 19014 6644 19066
rect 6668 19014 6698 19066
rect 6698 19014 6710 19066
rect 6710 19014 6724 19066
rect 6748 19014 6762 19066
rect 6762 19014 6774 19066
rect 6774 19014 6804 19066
rect 6828 19014 6838 19066
rect 6838 19014 6884 19066
rect 6588 19012 6644 19014
rect 6668 19012 6724 19014
rect 6748 19012 6804 19014
rect 6828 19012 6884 19014
rect 1398 2760 1454 2816
rect 2870 2080 2926 2136
rect 2962 1400 3018 1456
rect 2962 720 3018 776
rect 6588 17978 6644 17980
rect 6668 17978 6724 17980
rect 6748 17978 6804 17980
rect 6828 17978 6884 17980
rect 6588 17926 6634 17978
rect 6634 17926 6644 17978
rect 6668 17926 6698 17978
rect 6698 17926 6710 17978
rect 6710 17926 6724 17978
rect 6748 17926 6762 17978
rect 6762 17926 6774 17978
rect 6774 17926 6804 17978
rect 6828 17926 6838 17978
rect 6838 17926 6884 17978
rect 6588 17924 6644 17926
rect 6668 17924 6724 17926
rect 6748 17924 6804 17926
rect 6828 17924 6884 17926
rect 6588 16890 6644 16892
rect 6668 16890 6724 16892
rect 6748 16890 6804 16892
rect 6828 16890 6884 16892
rect 6588 16838 6634 16890
rect 6634 16838 6644 16890
rect 6668 16838 6698 16890
rect 6698 16838 6710 16890
rect 6710 16838 6724 16890
rect 6748 16838 6762 16890
rect 6762 16838 6774 16890
rect 6774 16838 6804 16890
rect 6828 16838 6838 16890
rect 6838 16838 6884 16890
rect 6588 16836 6644 16838
rect 6668 16836 6724 16838
rect 6748 16836 6804 16838
rect 6828 16836 6884 16838
rect 6588 15802 6644 15804
rect 6668 15802 6724 15804
rect 6748 15802 6804 15804
rect 6828 15802 6884 15804
rect 6588 15750 6634 15802
rect 6634 15750 6644 15802
rect 6668 15750 6698 15802
rect 6698 15750 6710 15802
rect 6710 15750 6724 15802
rect 6748 15750 6762 15802
rect 6762 15750 6774 15802
rect 6774 15750 6804 15802
rect 6828 15750 6838 15802
rect 6838 15750 6884 15802
rect 6588 15748 6644 15750
rect 6668 15748 6724 15750
rect 6748 15748 6804 15750
rect 6828 15748 6884 15750
rect 6588 14714 6644 14716
rect 6668 14714 6724 14716
rect 6748 14714 6804 14716
rect 6828 14714 6884 14716
rect 6588 14662 6634 14714
rect 6634 14662 6644 14714
rect 6668 14662 6698 14714
rect 6698 14662 6710 14714
rect 6710 14662 6724 14714
rect 6748 14662 6762 14714
rect 6762 14662 6774 14714
rect 6774 14662 6804 14714
rect 6828 14662 6838 14714
rect 6838 14662 6884 14714
rect 6588 14660 6644 14662
rect 6668 14660 6724 14662
rect 6748 14660 6804 14662
rect 6828 14660 6884 14662
rect 6588 13626 6644 13628
rect 6668 13626 6724 13628
rect 6748 13626 6804 13628
rect 6828 13626 6884 13628
rect 6588 13574 6634 13626
rect 6634 13574 6644 13626
rect 6668 13574 6698 13626
rect 6698 13574 6710 13626
rect 6710 13574 6724 13626
rect 6748 13574 6762 13626
rect 6762 13574 6774 13626
rect 6774 13574 6804 13626
rect 6828 13574 6838 13626
rect 6838 13574 6884 13626
rect 6588 13572 6644 13574
rect 6668 13572 6724 13574
rect 6748 13572 6804 13574
rect 6828 13572 6884 13574
rect 6588 12538 6644 12540
rect 6668 12538 6724 12540
rect 6748 12538 6804 12540
rect 6828 12538 6884 12540
rect 6588 12486 6634 12538
rect 6634 12486 6644 12538
rect 6668 12486 6698 12538
rect 6698 12486 6710 12538
rect 6710 12486 6724 12538
rect 6748 12486 6762 12538
rect 6762 12486 6774 12538
rect 6774 12486 6804 12538
rect 6828 12486 6838 12538
rect 6838 12486 6884 12538
rect 6588 12484 6644 12486
rect 6668 12484 6724 12486
rect 6748 12484 6804 12486
rect 6828 12484 6884 12486
rect 6588 11450 6644 11452
rect 6668 11450 6724 11452
rect 6748 11450 6804 11452
rect 6828 11450 6884 11452
rect 6588 11398 6634 11450
rect 6634 11398 6644 11450
rect 6668 11398 6698 11450
rect 6698 11398 6710 11450
rect 6710 11398 6724 11450
rect 6748 11398 6762 11450
rect 6762 11398 6774 11450
rect 6774 11398 6804 11450
rect 6828 11398 6838 11450
rect 6838 11398 6884 11450
rect 6588 11396 6644 11398
rect 6668 11396 6724 11398
rect 6748 11396 6804 11398
rect 6828 11396 6884 11398
rect 6588 10362 6644 10364
rect 6668 10362 6724 10364
rect 6748 10362 6804 10364
rect 6828 10362 6884 10364
rect 6588 10310 6634 10362
rect 6634 10310 6644 10362
rect 6668 10310 6698 10362
rect 6698 10310 6710 10362
rect 6710 10310 6724 10362
rect 6748 10310 6762 10362
rect 6762 10310 6774 10362
rect 6774 10310 6804 10362
rect 6828 10310 6838 10362
rect 6838 10310 6884 10362
rect 6588 10308 6644 10310
rect 6668 10308 6724 10310
rect 6748 10308 6804 10310
rect 6828 10308 6884 10310
rect 6588 9274 6644 9276
rect 6668 9274 6724 9276
rect 6748 9274 6804 9276
rect 6828 9274 6884 9276
rect 6588 9222 6634 9274
rect 6634 9222 6644 9274
rect 6668 9222 6698 9274
rect 6698 9222 6710 9274
rect 6710 9222 6724 9274
rect 6748 9222 6762 9274
rect 6762 9222 6774 9274
rect 6774 9222 6804 9274
rect 6828 9222 6838 9274
rect 6838 9222 6884 9274
rect 6588 9220 6644 9222
rect 6668 9220 6724 9222
rect 6748 9220 6804 9222
rect 6828 9220 6884 9222
rect 6588 8186 6644 8188
rect 6668 8186 6724 8188
rect 6748 8186 6804 8188
rect 6828 8186 6884 8188
rect 6588 8134 6634 8186
rect 6634 8134 6644 8186
rect 6668 8134 6698 8186
rect 6698 8134 6710 8186
rect 6710 8134 6724 8186
rect 6748 8134 6762 8186
rect 6762 8134 6774 8186
rect 6774 8134 6804 8186
rect 6828 8134 6838 8186
rect 6838 8134 6884 8186
rect 6588 8132 6644 8134
rect 6668 8132 6724 8134
rect 6748 8132 6804 8134
rect 6828 8132 6884 8134
rect 6588 7098 6644 7100
rect 6668 7098 6724 7100
rect 6748 7098 6804 7100
rect 6828 7098 6884 7100
rect 6588 7046 6634 7098
rect 6634 7046 6644 7098
rect 6668 7046 6698 7098
rect 6698 7046 6710 7098
rect 6710 7046 6724 7098
rect 6748 7046 6762 7098
rect 6762 7046 6774 7098
rect 6774 7046 6804 7098
rect 6828 7046 6838 7098
rect 6838 7046 6884 7098
rect 6588 7044 6644 7046
rect 6668 7044 6724 7046
rect 6748 7044 6804 7046
rect 6828 7044 6884 7046
rect 6588 6010 6644 6012
rect 6668 6010 6724 6012
rect 6748 6010 6804 6012
rect 6828 6010 6884 6012
rect 6588 5958 6634 6010
rect 6634 5958 6644 6010
rect 6668 5958 6698 6010
rect 6698 5958 6710 6010
rect 6710 5958 6724 6010
rect 6748 5958 6762 6010
rect 6762 5958 6774 6010
rect 6774 5958 6804 6010
rect 6828 5958 6838 6010
rect 6838 5958 6884 6010
rect 6588 5956 6644 5958
rect 6668 5956 6724 5958
rect 6748 5956 6804 5958
rect 6828 5956 6884 5958
rect 6588 4922 6644 4924
rect 6668 4922 6724 4924
rect 6748 4922 6804 4924
rect 6828 4922 6884 4924
rect 6588 4870 6634 4922
rect 6634 4870 6644 4922
rect 6668 4870 6698 4922
rect 6698 4870 6710 4922
rect 6710 4870 6724 4922
rect 6748 4870 6762 4922
rect 6762 4870 6774 4922
rect 6774 4870 6804 4922
rect 6828 4870 6838 4922
rect 6838 4870 6884 4922
rect 6588 4868 6644 4870
rect 6668 4868 6724 4870
rect 6748 4868 6804 4870
rect 6828 4868 6884 4870
rect 6588 3834 6644 3836
rect 6668 3834 6724 3836
rect 6748 3834 6804 3836
rect 6828 3834 6884 3836
rect 6588 3782 6634 3834
rect 6634 3782 6644 3834
rect 6668 3782 6698 3834
rect 6698 3782 6710 3834
rect 6710 3782 6724 3834
rect 6748 3782 6762 3834
rect 6762 3782 6774 3834
rect 6774 3782 6804 3834
rect 6828 3782 6838 3834
rect 6838 3782 6884 3834
rect 6588 3780 6644 3782
rect 6668 3780 6724 3782
rect 6748 3780 6804 3782
rect 6828 3780 6884 3782
rect 6588 2746 6644 2748
rect 6668 2746 6724 2748
rect 6748 2746 6804 2748
rect 6828 2746 6884 2748
rect 6588 2694 6634 2746
rect 6634 2694 6644 2746
rect 6668 2694 6698 2746
rect 6698 2694 6710 2746
rect 6710 2694 6724 2746
rect 6748 2694 6762 2746
rect 6762 2694 6774 2746
rect 6774 2694 6804 2746
rect 6828 2694 6838 2746
rect 6838 2694 6884 2746
rect 6588 2692 6644 2694
rect 6668 2692 6724 2694
rect 6748 2692 6804 2694
rect 6828 2692 6884 2694
rect 12220 33754 12276 33756
rect 12300 33754 12356 33756
rect 12380 33754 12436 33756
rect 12460 33754 12516 33756
rect 12220 33702 12266 33754
rect 12266 33702 12276 33754
rect 12300 33702 12330 33754
rect 12330 33702 12342 33754
rect 12342 33702 12356 33754
rect 12380 33702 12394 33754
rect 12394 33702 12406 33754
rect 12406 33702 12436 33754
rect 12460 33702 12470 33754
rect 12470 33702 12516 33754
rect 12220 33700 12276 33702
rect 12300 33700 12356 33702
rect 12380 33700 12436 33702
rect 12460 33700 12516 33702
rect 12220 32666 12276 32668
rect 12300 32666 12356 32668
rect 12380 32666 12436 32668
rect 12460 32666 12516 32668
rect 12220 32614 12266 32666
rect 12266 32614 12276 32666
rect 12300 32614 12330 32666
rect 12330 32614 12342 32666
rect 12342 32614 12356 32666
rect 12380 32614 12394 32666
rect 12394 32614 12406 32666
rect 12406 32614 12436 32666
rect 12460 32614 12470 32666
rect 12470 32614 12516 32666
rect 12220 32612 12276 32614
rect 12300 32612 12356 32614
rect 12380 32612 12436 32614
rect 12460 32612 12516 32614
rect 12220 31578 12276 31580
rect 12300 31578 12356 31580
rect 12380 31578 12436 31580
rect 12460 31578 12516 31580
rect 12220 31526 12266 31578
rect 12266 31526 12276 31578
rect 12300 31526 12330 31578
rect 12330 31526 12342 31578
rect 12342 31526 12356 31578
rect 12380 31526 12394 31578
rect 12394 31526 12406 31578
rect 12406 31526 12436 31578
rect 12460 31526 12470 31578
rect 12470 31526 12516 31578
rect 12220 31524 12276 31526
rect 12300 31524 12356 31526
rect 12380 31524 12436 31526
rect 12460 31524 12516 31526
rect 12220 30490 12276 30492
rect 12300 30490 12356 30492
rect 12380 30490 12436 30492
rect 12460 30490 12516 30492
rect 12220 30438 12266 30490
rect 12266 30438 12276 30490
rect 12300 30438 12330 30490
rect 12330 30438 12342 30490
rect 12342 30438 12356 30490
rect 12380 30438 12394 30490
rect 12394 30438 12406 30490
rect 12406 30438 12436 30490
rect 12460 30438 12470 30490
rect 12470 30438 12516 30490
rect 12220 30436 12276 30438
rect 12300 30436 12356 30438
rect 12380 30436 12436 30438
rect 12460 30436 12516 30438
rect 12220 29402 12276 29404
rect 12300 29402 12356 29404
rect 12380 29402 12436 29404
rect 12460 29402 12516 29404
rect 12220 29350 12266 29402
rect 12266 29350 12276 29402
rect 12300 29350 12330 29402
rect 12330 29350 12342 29402
rect 12342 29350 12356 29402
rect 12380 29350 12394 29402
rect 12394 29350 12406 29402
rect 12406 29350 12436 29402
rect 12460 29350 12470 29402
rect 12470 29350 12516 29402
rect 12220 29348 12276 29350
rect 12300 29348 12356 29350
rect 12380 29348 12436 29350
rect 12460 29348 12516 29350
rect 12220 28314 12276 28316
rect 12300 28314 12356 28316
rect 12380 28314 12436 28316
rect 12460 28314 12516 28316
rect 12220 28262 12266 28314
rect 12266 28262 12276 28314
rect 12300 28262 12330 28314
rect 12330 28262 12342 28314
rect 12342 28262 12356 28314
rect 12380 28262 12394 28314
rect 12394 28262 12406 28314
rect 12406 28262 12436 28314
rect 12460 28262 12470 28314
rect 12470 28262 12516 28314
rect 12220 28260 12276 28262
rect 12300 28260 12356 28262
rect 12380 28260 12436 28262
rect 12460 28260 12516 28262
rect 12220 27226 12276 27228
rect 12300 27226 12356 27228
rect 12380 27226 12436 27228
rect 12460 27226 12516 27228
rect 12220 27174 12266 27226
rect 12266 27174 12276 27226
rect 12300 27174 12330 27226
rect 12330 27174 12342 27226
rect 12342 27174 12356 27226
rect 12380 27174 12394 27226
rect 12394 27174 12406 27226
rect 12406 27174 12436 27226
rect 12460 27174 12470 27226
rect 12470 27174 12516 27226
rect 12220 27172 12276 27174
rect 12300 27172 12356 27174
rect 12380 27172 12436 27174
rect 12460 27172 12516 27174
rect 12220 26138 12276 26140
rect 12300 26138 12356 26140
rect 12380 26138 12436 26140
rect 12460 26138 12516 26140
rect 12220 26086 12266 26138
rect 12266 26086 12276 26138
rect 12300 26086 12330 26138
rect 12330 26086 12342 26138
rect 12342 26086 12356 26138
rect 12380 26086 12394 26138
rect 12394 26086 12406 26138
rect 12406 26086 12436 26138
rect 12460 26086 12470 26138
rect 12470 26086 12516 26138
rect 12220 26084 12276 26086
rect 12300 26084 12356 26086
rect 12380 26084 12436 26086
rect 12460 26084 12516 26086
rect 12220 25050 12276 25052
rect 12300 25050 12356 25052
rect 12380 25050 12436 25052
rect 12460 25050 12516 25052
rect 12220 24998 12266 25050
rect 12266 24998 12276 25050
rect 12300 24998 12330 25050
rect 12330 24998 12342 25050
rect 12342 24998 12356 25050
rect 12380 24998 12394 25050
rect 12394 24998 12406 25050
rect 12406 24998 12436 25050
rect 12460 24998 12470 25050
rect 12470 24998 12516 25050
rect 12220 24996 12276 24998
rect 12300 24996 12356 24998
rect 12380 24996 12436 24998
rect 12460 24996 12516 24998
rect 12220 23962 12276 23964
rect 12300 23962 12356 23964
rect 12380 23962 12436 23964
rect 12460 23962 12516 23964
rect 12220 23910 12266 23962
rect 12266 23910 12276 23962
rect 12300 23910 12330 23962
rect 12330 23910 12342 23962
rect 12342 23910 12356 23962
rect 12380 23910 12394 23962
rect 12394 23910 12406 23962
rect 12406 23910 12436 23962
rect 12460 23910 12470 23962
rect 12470 23910 12516 23962
rect 12220 23908 12276 23910
rect 12300 23908 12356 23910
rect 12380 23908 12436 23910
rect 12460 23908 12516 23910
rect 12220 22874 12276 22876
rect 12300 22874 12356 22876
rect 12380 22874 12436 22876
rect 12460 22874 12516 22876
rect 12220 22822 12266 22874
rect 12266 22822 12276 22874
rect 12300 22822 12330 22874
rect 12330 22822 12342 22874
rect 12342 22822 12356 22874
rect 12380 22822 12394 22874
rect 12394 22822 12406 22874
rect 12406 22822 12436 22874
rect 12460 22822 12470 22874
rect 12470 22822 12516 22874
rect 12220 22820 12276 22822
rect 12300 22820 12356 22822
rect 12380 22820 12436 22822
rect 12460 22820 12516 22822
rect 12220 21786 12276 21788
rect 12300 21786 12356 21788
rect 12380 21786 12436 21788
rect 12460 21786 12516 21788
rect 12220 21734 12266 21786
rect 12266 21734 12276 21786
rect 12300 21734 12330 21786
rect 12330 21734 12342 21786
rect 12342 21734 12356 21786
rect 12380 21734 12394 21786
rect 12394 21734 12406 21786
rect 12406 21734 12436 21786
rect 12460 21734 12470 21786
rect 12470 21734 12516 21786
rect 12220 21732 12276 21734
rect 12300 21732 12356 21734
rect 12380 21732 12436 21734
rect 12460 21732 12516 21734
rect 12220 20698 12276 20700
rect 12300 20698 12356 20700
rect 12380 20698 12436 20700
rect 12460 20698 12516 20700
rect 12220 20646 12266 20698
rect 12266 20646 12276 20698
rect 12300 20646 12330 20698
rect 12330 20646 12342 20698
rect 12342 20646 12356 20698
rect 12380 20646 12394 20698
rect 12394 20646 12406 20698
rect 12406 20646 12436 20698
rect 12460 20646 12470 20698
rect 12470 20646 12516 20698
rect 12220 20644 12276 20646
rect 12300 20644 12356 20646
rect 12380 20644 12436 20646
rect 12460 20644 12516 20646
rect 12220 19610 12276 19612
rect 12300 19610 12356 19612
rect 12380 19610 12436 19612
rect 12460 19610 12516 19612
rect 12220 19558 12266 19610
rect 12266 19558 12276 19610
rect 12300 19558 12330 19610
rect 12330 19558 12342 19610
rect 12342 19558 12356 19610
rect 12380 19558 12394 19610
rect 12394 19558 12406 19610
rect 12406 19558 12436 19610
rect 12460 19558 12470 19610
rect 12470 19558 12516 19610
rect 12220 19556 12276 19558
rect 12300 19556 12356 19558
rect 12380 19556 12436 19558
rect 12460 19556 12516 19558
rect 12220 18522 12276 18524
rect 12300 18522 12356 18524
rect 12380 18522 12436 18524
rect 12460 18522 12516 18524
rect 12220 18470 12266 18522
rect 12266 18470 12276 18522
rect 12300 18470 12330 18522
rect 12330 18470 12342 18522
rect 12342 18470 12356 18522
rect 12380 18470 12394 18522
rect 12394 18470 12406 18522
rect 12406 18470 12436 18522
rect 12460 18470 12470 18522
rect 12470 18470 12516 18522
rect 12220 18468 12276 18470
rect 12300 18468 12356 18470
rect 12380 18468 12436 18470
rect 12460 18468 12516 18470
rect 15290 31864 15346 31920
rect 12220 17434 12276 17436
rect 12300 17434 12356 17436
rect 12380 17434 12436 17436
rect 12460 17434 12516 17436
rect 12220 17382 12266 17434
rect 12266 17382 12276 17434
rect 12300 17382 12330 17434
rect 12330 17382 12342 17434
rect 12342 17382 12356 17434
rect 12380 17382 12394 17434
rect 12394 17382 12406 17434
rect 12406 17382 12436 17434
rect 12460 17382 12470 17434
rect 12470 17382 12516 17434
rect 12220 17380 12276 17382
rect 12300 17380 12356 17382
rect 12380 17380 12436 17382
rect 12460 17380 12516 17382
rect 12220 16346 12276 16348
rect 12300 16346 12356 16348
rect 12380 16346 12436 16348
rect 12460 16346 12516 16348
rect 12220 16294 12266 16346
rect 12266 16294 12276 16346
rect 12300 16294 12330 16346
rect 12330 16294 12342 16346
rect 12342 16294 12356 16346
rect 12380 16294 12394 16346
rect 12394 16294 12406 16346
rect 12406 16294 12436 16346
rect 12460 16294 12470 16346
rect 12470 16294 12516 16346
rect 12220 16292 12276 16294
rect 12300 16292 12356 16294
rect 12380 16292 12436 16294
rect 12460 16292 12516 16294
rect 12220 15258 12276 15260
rect 12300 15258 12356 15260
rect 12380 15258 12436 15260
rect 12460 15258 12516 15260
rect 12220 15206 12266 15258
rect 12266 15206 12276 15258
rect 12300 15206 12330 15258
rect 12330 15206 12342 15258
rect 12342 15206 12356 15258
rect 12380 15206 12394 15258
rect 12394 15206 12406 15258
rect 12406 15206 12436 15258
rect 12460 15206 12470 15258
rect 12470 15206 12516 15258
rect 12220 15204 12276 15206
rect 12300 15204 12356 15206
rect 12380 15204 12436 15206
rect 12460 15204 12516 15206
rect 12220 14170 12276 14172
rect 12300 14170 12356 14172
rect 12380 14170 12436 14172
rect 12460 14170 12516 14172
rect 12220 14118 12266 14170
rect 12266 14118 12276 14170
rect 12300 14118 12330 14170
rect 12330 14118 12342 14170
rect 12342 14118 12356 14170
rect 12380 14118 12394 14170
rect 12394 14118 12406 14170
rect 12406 14118 12436 14170
rect 12460 14118 12470 14170
rect 12470 14118 12516 14170
rect 12220 14116 12276 14118
rect 12300 14116 12356 14118
rect 12380 14116 12436 14118
rect 12460 14116 12516 14118
rect 12220 13082 12276 13084
rect 12300 13082 12356 13084
rect 12380 13082 12436 13084
rect 12460 13082 12516 13084
rect 12220 13030 12266 13082
rect 12266 13030 12276 13082
rect 12300 13030 12330 13082
rect 12330 13030 12342 13082
rect 12342 13030 12356 13082
rect 12380 13030 12394 13082
rect 12394 13030 12406 13082
rect 12406 13030 12436 13082
rect 12460 13030 12470 13082
rect 12470 13030 12516 13082
rect 12220 13028 12276 13030
rect 12300 13028 12356 13030
rect 12380 13028 12436 13030
rect 12460 13028 12516 13030
rect 12220 11994 12276 11996
rect 12300 11994 12356 11996
rect 12380 11994 12436 11996
rect 12460 11994 12516 11996
rect 12220 11942 12266 11994
rect 12266 11942 12276 11994
rect 12300 11942 12330 11994
rect 12330 11942 12342 11994
rect 12342 11942 12356 11994
rect 12380 11942 12394 11994
rect 12394 11942 12406 11994
rect 12406 11942 12436 11994
rect 12460 11942 12470 11994
rect 12470 11942 12516 11994
rect 12220 11940 12276 11942
rect 12300 11940 12356 11942
rect 12380 11940 12436 11942
rect 12460 11940 12516 11942
rect 12220 10906 12276 10908
rect 12300 10906 12356 10908
rect 12380 10906 12436 10908
rect 12460 10906 12516 10908
rect 12220 10854 12266 10906
rect 12266 10854 12276 10906
rect 12300 10854 12330 10906
rect 12330 10854 12342 10906
rect 12342 10854 12356 10906
rect 12380 10854 12394 10906
rect 12394 10854 12406 10906
rect 12406 10854 12436 10906
rect 12460 10854 12470 10906
rect 12470 10854 12516 10906
rect 12220 10852 12276 10854
rect 12300 10852 12356 10854
rect 12380 10852 12436 10854
rect 12460 10852 12516 10854
rect 12220 9818 12276 9820
rect 12300 9818 12356 9820
rect 12380 9818 12436 9820
rect 12460 9818 12516 9820
rect 12220 9766 12266 9818
rect 12266 9766 12276 9818
rect 12300 9766 12330 9818
rect 12330 9766 12342 9818
rect 12342 9766 12356 9818
rect 12380 9766 12394 9818
rect 12394 9766 12406 9818
rect 12406 9766 12436 9818
rect 12460 9766 12470 9818
rect 12470 9766 12516 9818
rect 12220 9764 12276 9766
rect 12300 9764 12356 9766
rect 12380 9764 12436 9766
rect 12460 9764 12516 9766
rect 12220 8730 12276 8732
rect 12300 8730 12356 8732
rect 12380 8730 12436 8732
rect 12460 8730 12516 8732
rect 12220 8678 12266 8730
rect 12266 8678 12276 8730
rect 12300 8678 12330 8730
rect 12330 8678 12342 8730
rect 12342 8678 12356 8730
rect 12380 8678 12394 8730
rect 12394 8678 12406 8730
rect 12406 8678 12436 8730
rect 12460 8678 12470 8730
rect 12470 8678 12516 8730
rect 12220 8676 12276 8678
rect 12300 8676 12356 8678
rect 12380 8676 12436 8678
rect 12460 8676 12516 8678
rect 12220 7642 12276 7644
rect 12300 7642 12356 7644
rect 12380 7642 12436 7644
rect 12460 7642 12516 7644
rect 12220 7590 12266 7642
rect 12266 7590 12276 7642
rect 12300 7590 12330 7642
rect 12330 7590 12342 7642
rect 12342 7590 12356 7642
rect 12380 7590 12394 7642
rect 12394 7590 12406 7642
rect 12406 7590 12436 7642
rect 12460 7590 12470 7642
rect 12470 7590 12516 7642
rect 12220 7588 12276 7590
rect 12300 7588 12356 7590
rect 12380 7588 12436 7590
rect 12460 7588 12516 7590
rect 12220 6554 12276 6556
rect 12300 6554 12356 6556
rect 12380 6554 12436 6556
rect 12460 6554 12516 6556
rect 12220 6502 12266 6554
rect 12266 6502 12276 6554
rect 12300 6502 12330 6554
rect 12330 6502 12342 6554
rect 12342 6502 12356 6554
rect 12380 6502 12394 6554
rect 12394 6502 12406 6554
rect 12406 6502 12436 6554
rect 12460 6502 12470 6554
rect 12470 6502 12516 6554
rect 12220 6500 12276 6502
rect 12300 6500 12356 6502
rect 12380 6500 12436 6502
rect 12460 6500 12516 6502
rect 12220 5466 12276 5468
rect 12300 5466 12356 5468
rect 12380 5466 12436 5468
rect 12460 5466 12516 5468
rect 12220 5414 12266 5466
rect 12266 5414 12276 5466
rect 12300 5414 12330 5466
rect 12330 5414 12342 5466
rect 12342 5414 12356 5466
rect 12380 5414 12394 5466
rect 12394 5414 12406 5466
rect 12406 5414 12436 5466
rect 12460 5414 12470 5466
rect 12470 5414 12516 5466
rect 12220 5412 12276 5414
rect 12300 5412 12356 5414
rect 12380 5412 12436 5414
rect 12460 5412 12516 5414
rect 12220 4378 12276 4380
rect 12300 4378 12356 4380
rect 12380 4378 12436 4380
rect 12460 4378 12516 4380
rect 12220 4326 12266 4378
rect 12266 4326 12276 4378
rect 12300 4326 12330 4378
rect 12330 4326 12342 4378
rect 12342 4326 12356 4378
rect 12380 4326 12394 4378
rect 12394 4326 12406 4378
rect 12406 4326 12436 4378
rect 12460 4326 12470 4378
rect 12470 4326 12516 4378
rect 12220 4324 12276 4326
rect 12300 4324 12356 4326
rect 12380 4324 12436 4326
rect 12460 4324 12516 4326
rect 12220 3290 12276 3292
rect 12300 3290 12356 3292
rect 12380 3290 12436 3292
rect 12460 3290 12516 3292
rect 12220 3238 12266 3290
rect 12266 3238 12276 3290
rect 12300 3238 12330 3290
rect 12330 3238 12342 3290
rect 12342 3238 12356 3290
rect 12380 3238 12394 3290
rect 12394 3238 12406 3290
rect 12406 3238 12436 3290
rect 12460 3238 12470 3290
rect 12470 3238 12516 3290
rect 12220 3236 12276 3238
rect 12300 3236 12356 3238
rect 12380 3236 12436 3238
rect 12460 3236 12516 3238
rect 12220 2202 12276 2204
rect 12300 2202 12356 2204
rect 12380 2202 12436 2204
rect 12460 2202 12516 2204
rect 12220 2150 12266 2202
rect 12266 2150 12276 2202
rect 12300 2150 12330 2202
rect 12330 2150 12342 2202
rect 12342 2150 12356 2202
rect 12380 2150 12394 2202
rect 12394 2150 12406 2202
rect 12406 2150 12436 2202
rect 12460 2150 12470 2202
rect 12470 2150 12516 2202
rect 12220 2148 12276 2150
rect 12300 2148 12356 2150
rect 12380 2148 12436 2150
rect 12460 2148 12516 2150
rect 17852 33210 17908 33212
rect 17932 33210 17988 33212
rect 18012 33210 18068 33212
rect 18092 33210 18148 33212
rect 17852 33158 17898 33210
rect 17898 33158 17908 33210
rect 17932 33158 17962 33210
rect 17962 33158 17974 33210
rect 17974 33158 17988 33210
rect 18012 33158 18026 33210
rect 18026 33158 18038 33210
rect 18038 33158 18068 33210
rect 18092 33158 18102 33210
rect 18102 33158 18148 33210
rect 17852 33156 17908 33158
rect 17932 33156 17988 33158
rect 18012 33156 18068 33158
rect 18092 33156 18148 33158
rect 17852 32122 17908 32124
rect 17932 32122 17988 32124
rect 18012 32122 18068 32124
rect 18092 32122 18148 32124
rect 17852 32070 17898 32122
rect 17898 32070 17908 32122
rect 17932 32070 17962 32122
rect 17962 32070 17974 32122
rect 17974 32070 17988 32122
rect 18012 32070 18026 32122
rect 18026 32070 18038 32122
rect 18038 32070 18068 32122
rect 18092 32070 18102 32122
rect 18102 32070 18148 32122
rect 17852 32068 17908 32070
rect 17932 32068 17988 32070
rect 18012 32068 18068 32070
rect 18092 32068 18148 32070
rect 17852 31034 17908 31036
rect 17932 31034 17988 31036
rect 18012 31034 18068 31036
rect 18092 31034 18148 31036
rect 17852 30982 17898 31034
rect 17898 30982 17908 31034
rect 17932 30982 17962 31034
rect 17962 30982 17974 31034
rect 17974 30982 17988 31034
rect 18012 30982 18026 31034
rect 18026 30982 18038 31034
rect 18038 30982 18068 31034
rect 18092 30982 18102 31034
rect 18102 30982 18148 31034
rect 17852 30980 17908 30982
rect 17932 30980 17988 30982
rect 18012 30980 18068 30982
rect 18092 30980 18148 30982
rect 17852 29946 17908 29948
rect 17932 29946 17988 29948
rect 18012 29946 18068 29948
rect 18092 29946 18148 29948
rect 17852 29894 17898 29946
rect 17898 29894 17908 29946
rect 17932 29894 17962 29946
rect 17962 29894 17974 29946
rect 17974 29894 17988 29946
rect 18012 29894 18026 29946
rect 18026 29894 18038 29946
rect 18038 29894 18068 29946
rect 18092 29894 18102 29946
rect 18102 29894 18148 29946
rect 17852 29892 17908 29894
rect 17932 29892 17988 29894
rect 18012 29892 18068 29894
rect 18092 29892 18148 29894
rect 17852 28858 17908 28860
rect 17932 28858 17988 28860
rect 18012 28858 18068 28860
rect 18092 28858 18148 28860
rect 17852 28806 17898 28858
rect 17898 28806 17908 28858
rect 17932 28806 17962 28858
rect 17962 28806 17974 28858
rect 17974 28806 17988 28858
rect 18012 28806 18026 28858
rect 18026 28806 18038 28858
rect 18038 28806 18068 28858
rect 18092 28806 18102 28858
rect 18102 28806 18148 28858
rect 17852 28804 17908 28806
rect 17932 28804 17988 28806
rect 18012 28804 18068 28806
rect 18092 28804 18148 28806
rect 17852 27770 17908 27772
rect 17932 27770 17988 27772
rect 18012 27770 18068 27772
rect 18092 27770 18148 27772
rect 17852 27718 17898 27770
rect 17898 27718 17908 27770
rect 17932 27718 17962 27770
rect 17962 27718 17974 27770
rect 17974 27718 17988 27770
rect 18012 27718 18026 27770
rect 18026 27718 18038 27770
rect 18038 27718 18068 27770
rect 18092 27718 18102 27770
rect 18102 27718 18148 27770
rect 17852 27716 17908 27718
rect 17932 27716 17988 27718
rect 18012 27716 18068 27718
rect 18092 27716 18148 27718
rect 17852 26682 17908 26684
rect 17932 26682 17988 26684
rect 18012 26682 18068 26684
rect 18092 26682 18148 26684
rect 17852 26630 17898 26682
rect 17898 26630 17908 26682
rect 17932 26630 17962 26682
rect 17962 26630 17974 26682
rect 17974 26630 17988 26682
rect 18012 26630 18026 26682
rect 18026 26630 18038 26682
rect 18038 26630 18068 26682
rect 18092 26630 18102 26682
rect 18102 26630 18148 26682
rect 17852 26628 17908 26630
rect 17932 26628 17988 26630
rect 18012 26628 18068 26630
rect 18092 26628 18148 26630
rect 17852 25594 17908 25596
rect 17932 25594 17988 25596
rect 18012 25594 18068 25596
rect 18092 25594 18148 25596
rect 17852 25542 17898 25594
rect 17898 25542 17908 25594
rect 17932 25542 17962 25594
rect 17962 25542 17974 25594
rect 17974 25542 17988 25594
rect 18012 25542 18026 25594
rect 18026 25542 18038 25594
rect 18038 25542 18068 25594
rect 18092 25542 18102 25594
rect 18102 25542 18148 25594
rect 17852 25540 17908 25542
rect 17932 25540 17988 25542
rect 18012 25540 18068 25542
rect 18092 25540 18148 25542
rect 17852 24506 17908 24508
rect 17932 24506 17988 24508
rect 18012 24506 18068 24508
rect 18092 24506 18148 24508
rect 17852 24454 17898 24506
rect 17898 24454 17908 24506
rect 17932 24454 17962 24506
rect 17962 24454 17974 24506
rect 17974 24454 17988 24506
rect 18012 24454 18026 24506
rect 18026 24454 18038 24506
rect 18038 24454 18068 24506
rect 18092 24454 18102 24506
rect 18102 24454 18148 24506
rect 17852 24452 17908 24454
rect 17932 24452 17988 24454
rect 18012 24452 18068 24454
rect 18092 24452 18148 24454
rect 17852 23418 17908 23420
rect 17932 23418 17988 23420
rect 18012 23418 18068 23420
rect 18092 23418 18148 23420
rect 17852 23366 17898 23418
rect 17898 23366 17908 23418
rect 17932 23366 17962 23418
rect 17962 23366 17974 23418
rect 17974 23366 17988 23418
rect 18012 23366 18026 23418
rect 18026 23366 18038 23418
rect 18038 23366 18068 23418
rect 18092 23366 18102 23418
rect 18102 23366 18148 23418
rect 17852 23364 17908 23366
rect 17932 23364 17988 23366
rect 18012 23364 18068 23366
rect 18092 23364 18148 23366
rect 17852 22330 17908 22332
rect 17932 22330 17988 22332
rect 18012 22330 18068 22332
rect 18092 22330 18148 22332
rect 17852 22278 17898 22330
rect 17898 22278 17908 22330
rect 17932 22278 17962 22330
rect 17962 22278 17974 22330
rect 17974 22278 17988 22330
rect 18012 22278 18026 22330
rect 18026 22278 18038 22330
rect 18038 22278 18068 22330
rect 18092 22278 18102 22330
rect 18102 22278 18148 22330
rect 17852 22276 17908 22278
rect 17932 22276 17988 22278
rect 18012 22276 18068 22278
rect 18092 22276 18148 22278
rect 17852 21242 17908 21244
rect 17932 21242 17988 21244
rect 18012 21242 18068 21244
rect 18092 21242 18148 21244
rect 17852 21190 17898 21242
rect 17898 21190 17908 21242
rect 17932 21190 17962 21242
rect 17962 21190 17974 21242
rect 17974 21190 17988 21242
rect 18012 21190 18026 21242
rect 18026 21190 18038 21242
rect 18038 21190 18068 21242
rect 18092 21190 18102 21242
rect 18102 21190 18148 21242
rect 17852 21188 17908 21190
rect 17932 21188 17988 21190
rect 18012 21188 18068 21190
rect 18092 21188 18148 21190
rect 17852 20154 17908 20156
rect 17932 20154 17988 20156
rect 18012 20154 18068 20156
rect 18092 20154 18148 20156
rect 17852 20102 17898 20154
rect 17898 20102 17908 20154
rect 17932 20102 17962 20154
rect 17962 20102 17974 20154
rect 17974 20102 17988 20154
rect 18012 20102 18026 20154
rect 18026 20102 18038 20154
rect 18038 20102 18068 20154
rect 18092 20102 18102 20154
rect 18102 20102 18148 20154
rect 17852 20100 17908 20102
rect 17932 20100 17988 20102
rect 18012 20100 18068 20102
rect 18092 20100 18148 20102
rect 17852 19066 17908 19068
rect 17932 19066 17988 19068
rect 18012 19066 18068 19068
rect 18092 19066 18148 19068
rect 17852 19014 17898 19066
rect 17898 19014 17908 19066
rect 17932 19014 17962 19066
rect 17962 19014 17974 19066
rect 17974 19014 17988 19066
rect 18012 19014 18026 19066
rect 18026 19014 18038 19066
rect 18038 19014 18068 19066
rect 18092 19014 18102 19066
rect 18102 19014 18148 19066
rect 17852 19012 17908 19014
rect 17932 19012 17988 19014
rect 18012 19012 18068 19014
rect 18092 19012 18148 19014
rect 17852 17978 17908 17980
rect 17932 17978 17988 17980
rect 18012 17978 18068 17980
rect 18092 17978 18148 17980
rect 17852 17926 17898 17978
rect 17898 17926 17908 17978
rect 17932 17926 17962 17978
rect 17962 17926 17974 17978
rect 17974 17926 17988 17978
rect 18012 17926 18026 17978
rect 18026 17926 18038 17978
rect 18038 17926 18068 17978
rect 18092 17926 18102 17978
rect 18102 17926 18148 17978
rect 17852 17924 17908 17926
rect 17932 17924 17988 17926
rect 18012 17924 18068 17926
rect 18092 17924 18148 17926
rect 17852 16890 17908 16892
rect 17932 16890 17988 16892
rect 18012 16890 18068 16892
rect 18092 16890 18148 16892
rect 17852 16838 17898 16890
rect 17898 16838 17908 16890
rect 17932 16838 17962 16890
rect 17962 16838 17974 16890
rect 17974 16838 17988 16890
rect 18012 16838 18026 16890
rect 18026 16838 18038 16890
rect 18038 16838 18068 16890
rect 18092 16838 18102 16890
rect 18102 16838 18148 16890
rect 17852 16836 17908 16838
rect 17932 16836 17988 16838
rect 18012 16836 18068 16838
rect 18092 16836 18148 16838
rect 17852 15802 17908 15804
rect 17932 15802 17988 15804
rect 18012 15802 18068 15804
rect 18092 15802 18148 15804
rect 17852 15750 17898 15802
rect 17898 15750 17908 15802
rect 17932 15750 17962 15802
rect 17962 15750 17974 15802
rect 17974 15750 17988 15802
rect 18012 15750 18026 15802
rect 18026 15750 18038 15802
rect 18038 15750 18068 15802
rect 18092 15750 18102 15802
rect 18102 15750 18148 15802
rect 17852 15748 17908 15750
rect 17932 15748 17988 15750
rect 18012 15748 18068 15750
rect 18092 15748 18148 15750
rect 17852 14714 17908 14716
rect 17932 14714 17988 14716
rect 18012 14714 18068 14716
rect 18092 14714 18148 14716
rect 17852 14662 17898 14714
rect 17898 14662 17908 14714
rect 17932 14662 17962 14714
rect 17962 14662 17974 14714
rect 17974 14662 17988 14714
rect 18012 14662 18026 14714
rect 18026 14662 18038 14714
rect 18038 14662 18068 14714
rect 18092 14662 18102 14714
rect 18102 14662 18148 14714
rect 17852 14660 17908 14662
rect 17932 14660 17988 14662
rect 18012 14660 18068 14662
rect 18092 14660 18148 14662
rect 17852 13626 17908 13628
rect 17932 13626 17988 13628
rect 18012 13626 18068 13628
rect 18092 13626 18148 13628
rect 17852 13574 17898 13626
rect 17898 13574 17908 13626
rect 17932 13574 17962 13626
rect 17962 13574 17974 13626
rect 17974 13574 17988 13626
rect 18012 13574 18026 13626
rect 18026 13574 18038 13626
rect 18038 13574 18068 13626
rect 18092 13574 18102 13626
rect 18102 13574 18148 13626
rect 17852 13572 17908 13574
rect 17932 13572 17988 13574
rect 18012 13572 18068 13574
rect 18092 13572 18148 13574
rect 17852 12538 17908 12540
rect 17932 12538 17988 12540
rect 18012 12538 18068 12540
rect 18092 12538 18148 12540
rect 17852 12486 17898 12538
rect 17898 12486 17908 12538
rect 17932 12486 17962 12538
rect 17962 12486 17974 12538
rect 17974 12486 17988 12538
rect 18012 12486 18026 12538
rect 18026 12486 18038 12538
rect 18038 12486 18068 12538
rect 18092 12486 18102 12538
rect 18102 12486 18148 12538
rect 17852 12484 17908 12486
rect 17932 12484 17988 12486
rect 18012 12484 18068 12486
rect 18092 12484 18148 12486
rect 17852 11450 17908 11452
rect 17932 11450 17988 11452
rect 18012 11450 18068 11452
rect 18092 11450 18148 11452
rect 17852 11398 17898 11450
rect 17898 11398 17908 11450
rect 17932 11398 17962 11450
rect 17962 11398 17974 11450
rect 17974 11398 17988 11450
rect 18012 11398 18026 11450
rect 18026 11398 18038 11450
rect 18038 11398 18068 11450
rect 18092 11398 18102 11450
rect 18102 11398 18148 11450
rect 17852 11396 17908 11398
rect 17932 11396 17988 11398
rect 18012 11396 18068 11398
rect 18092 11396 18148 11398
rect 17852 10362 17908 10364
rect 17932 10362 17988 10364
rect 18012 10362 18068 10364
rect 18092 10362 18148 10364
rect 17852 10310 17898 10362
rect 17898 10310 17908 10362
rect 17932 10310 17962 10362
rect 17962 10310 17974 10362
rect 17974 10310 17988 10362
rect 18012 10310 18026 10362
rect 18026 10310 18038 10362
rect 18038 10310 18068 10362
rect 18092 10310 18102 10362
rect 18102 10310 18148 10362
rect 17852 10308 17908 10310
rect 17932 10308 17988 10310
rect 18012 10308 18068 10310
rect 18092 10308 18148 10310
rect 17852 9274 17908 9276
rect 17932 9274 17988 9276
rect 18012 9274 18068 9276
rect 18092 9274 18148 9276
rect 17852 9222 17898 9274
rect 17898 9222 17908 9274
rect 17932 9222 17962 9274
rect 17962 9222 17974 9274
rect 17974 9222 17988 9274
rect 18012 9222 18026 9274
rect 18026 9222 18038 9274
rect 18038 9222 18068 9274
rect 18092 9222 18102 9274
rect 18102 9222 18148 9274
rect 17852 9220 17908 9222
rect 17932 9220 17988 9222
rect 18012 9220 18068 9222
rect 18092 9220 18148 9222
rect 17852 8186 17908 8188
rect 17932 8186 17988 8188
rect 18012 8186 18068 8188
rect 18092 8186 18148 8188
rect 17852 8134 17898 8186
rect 17898 8134 17908 8186
rect 17932 8134 17962 8186
rect 17962 8134 17974 8186
rect 17974 8134 17988 8186
rect 18012 8134 18026 8186
rect 18026 8134 18038 8186
rect 18038 8134 18068 8186
rect 18092 8134 18102 8186
rect 18102 8134 18148 8186
rect 17852 8132 17908 8134
rect 17932 8132 17988 8134
rect 18012 8132 18068 8134
rect 18092 8132 18148 8134
rect 17852 7098 17908 7100
rect 17932 7098 17988 7100
rect 18012 7098 18068 7100
rect 18092 7098 18148 7100
rect 17852 7046 17898 7098
rect 17898 7046 17908 7098
rect 17932 7046 17962 7098
rect 17962 7046 17974 7098
rect 17974 7046 17988 7098
rect 18012 7046 18026 7098
rect 18026 7046 18038 7098
rect 18038 7046 18068 7098
rect 18092 7046 18102 7098
rect 18102 7046 18148 7098
rect 17852 7044 17908 7046
rect 17932 7044 17988 7046
rect 18012 7044 18068 7046
rect 18092 7044 18148 7046
rect 17852 6010 17908 6012
rect 17932 6010 17988 6012
rect 18012 6010 18068 6012
rect 18092 6010 18148 6012
rect 17852 5958 17898 6010
rect 17898 5958 17908 6010
rect 17932 5958 17962 6010
rect 17962 5958 17974 6010
rect 17974 5958 17988 6010
rect 18012 5958 18026 6010
rect 18026 5958 18038 6010
rect 18038 5958 18068 6010
rect 18092 5958 18102 6010
rect 18102 5958 18148 6010
rect 17852 5956 17908 5958
rect 17932 5956 17988 5958
rect 18012 5956 18068 5958
rect 18092 5956 18148 5958
rect 17852 4922 17908 4924
rect 17932 4922 17988 4924
rect 18012 4922 18068 4924
rect 18092 4922 18148 4924
rect 17852 4870 17898 4922
rect 17898 4870 17908 4922
rect 17932 4870 17962 4922
rect 17962 4870 17974 4922
rect 17974 4870 17988 4922
rect 18012 4870 18026 4922
rect 18026 4870 18038 4922
rect 18038 4870 18068 4922
rect 18092 4870 18102 4922
rect 18102 4870 18148 4922
rect 17852 4868 17908 4870
rect 17932 4868 17988 4870
rect 18012 4868 18068 4870
rect 18092 4868 18148 4870
rect 17852 3834 17908 3836
rect 17932 3834 17988 3836
rect 18012 3834 18068 3836
rect 18092 3834 18148 3836
rect 17852 3782 17898 3834
rect 17898 3782 17908 3834
rect 17932 3782 17962 3834
rect 17962 3782 17974 3834
rect 17974 3782 17988 3834
rect 18012 3782 18026 3834
rect 18026 3782 18038 3834
rect 18038 3782 18068 3834
rect 18092 3782 18102 3834
rect 18102 3782 18148 3834
rect 17852 3780 17908 3782
rect 17932 3780 17988 3782
rect 18012 3780 18068 3782
rect 18092 3780 18148 3782
rect 17852 2746 17908 2748
rect 17932 2746 17988 2748
rect 18012 2746 18068 2748
rect 18092 2746 18148 2748
rect 17852 2694 17898 2746
rect 17898 2694 17908 2746
rect 17932 2694 17962 2746
rect 17962 2694 17974 2746
rect 17974 2694 17988 2746
rect 18012 2694 18026 2746
rect 18026 2694 18038 2746
rect 18038 2694 18068 2746
rect 18092 2694 18102 2746
rect 18102 2694 18148 2746
rect 17852 2692 17908 2694
rect 17932 2692 17988 2694
rect 18012 2692 18068 2694
rect 18092 2692 18148 2694
rect 19062 3440 19118 3496
rect 23484 33754 23540 33756
rect 23564 33754 23620 33756
rect 23644 33754 23700 33756
rect 23724 33754 23780 33756
rect 23484 33702 23530 33754
rect 23530 33702 23540 33754
rect 23564 33702 23594 33754
rect 23594 33702 23606 33754
rect 23606 33702 23620 33754
rect 23644 33702 23658 33754
rect 23658 33702 23670 33754
rect 23670 33702 23700 33754
rect 23724 33702 23734 33754
rect 23734 33702 23780 33754
rect 23484 33700 23540 33702
rect 23564 33700 23620 33702
rect 23644 33700 23700 33702
rect 23724 33700 23780 33702
rect 23484 32666 23540 32668
rect 23564 32666 23620 32668
rect 23644 32666 23700 32668
rect 23724 32666 23780 32668
rect 23484 32614 23530 32666
rect 23530 32614 23540 32666
rect 23564 32614 23594 32666
rect 23594 32614 23606 32666
rect 23606 32614 23620 32666
rect 23644 32614 23658 32666
rect 23658 32614 23670 32666
rect 23670 32614 23700 32666
rect 23724 32614 23734 32666
rect 23734 32614 23780 32666
rect 23484 32612 23540 32614
rect 23564 32612 23620 32614
rect 23644 32612 23700 32614
rect 23724 32612 23780 32614
rect 23484 31578 23540 31580
rect 23564 31578 23620 31580
rect 23644 31578 23700 31580
rect 23724 31578 23780 31580
rect 23484 31526 23530 31578
rect 23530 31526 23540 31578
rect 23564 31526 23594 31578
rect 23594 31526 23606 31578
rect 23606 31526 23620 31578
rect 23644 31526 23658 31578
rect 23658 31526 23670 31578
rect 23670 31526 23700 31578
rect 23724 31526 23734 31578
rect 23734 31526 23780 31578
rect 23484 31524 23540 31526
rect 23564 31524 23620 31526
rect 23644 31524 23700 31526
rect 23724 31524 23780 31526
rect 23484 30490 23540 30492
rect 23564 30490 23620 30492
rect 23644 30490 23700 30492
rect 23724 30490 23780 30492
rect 23484 30438 23530 30490
rect 23530 30438 23540 30490
rect 23564 30438 23594 30490
rect 23594 30438 23606 30490
rect 23606 30438 23620 30490
rect 23644 30438 23658 30490
rect 23658 30438 23670 30490
rect 23670 30438 23700 30490
rect 23724 30438 23734 30490
rect 23734 30438 23780 30490
rect 23484 30436 23540 30438
rect 23564 30436 23620 30438
rect 23644 30436 23700 30438
rect 23724 30436 23780 30438
rect 23484 29402 23540 29404
rect 23564 29402 23620 29404
rect 23644 29402 23700 29404
rect 23724 29402 23780 29404
rect 23484 29350 23530 29402
rect 23530 29350 23540 29402
rect 23564 29350 23594 29402
rect 23594 29350 23606 29402
rect 23606 29350 23620 29402
rect 23644 29350 23658 29402
rect 23658 29350 23670 29402
rect 23670 29350 23700 29402
rect 23724 29350 23734 29402
rect 23734 29350 23780 29402
rect 23484 29348 23540 29350
rect 23564 29348 23620 29350
rect 23644 29348 23700 29350
rect 23724 29348 23780 29350
rect 23484 28314 23540 28316
rect 23564 28314 23620 28316
rect 23644 28314 23700 28316
rect 23724 28314 23780 28316
rect 23484 28262 23530 28314
rect 23530 28262 23540 28314
rect 23564 28262 23594 28314
rect 23594 28262 23606 28314
rect 23606 28262 23620 28314
rect 23644 28262 23658 28314
rect 23658 28262 23670 28314
rect 23670 28262 23700 28314
rect 23724 28262 23734 28314
rect 23734 28262 23780 28314
rect 23484 28260 23540 28262
rect 23564 28260 23620 28262
rect 23644 28260 23700 28262
rect 23724 28260 23780 28262
rect 23484 27226 23540 27228
rect 23564 27226 23620 27228
rect 23644 27226 23700 27228
rect 23724 27226 23780 27228
rect 23484 27174 23530 27226
rect 23530 27174 23540 27226
rect 23564 27174 23594 27226
rect 23594 27174 23606 27226
rect 23606 27174 23620 27226
rect 23644 27174 23658 27226
rect 23658 27174 23670 27226
rect 23670 27174 23700 27226
rect 23724 27174 23734 27226
rect 23734 27174 23780 27226
rect 23484 27172 23540 27174
rect 23564 27172 23620 27174
rect 23644 27172 23700 27174
rect 23724 27172 23780 27174
rect 23484 26138 23540 26140
rect 23564 26138 23620 26140
rect 23644 26138 23700 26140
rect 23724 26138 23780 26140
rect 23484 26086 23530 26138
rect 23530 26086 23540 26138
rect 23564 26086 23594 26138
rect 23594 26086 23606 26138
rect 23606 26086 23620 26138
rect 23644 26086 23658 26138
rect 23658 26086 23670 26138
rect 23670 26086 23700 26138
rect 23724 26086 23734 26138
rect 23734 26086 23780 26138
rect 23484 26084 23540 26086
rect 23564 26084 23620 26086
rect 23644 26084 23700 26086
rect 23724 26084 23780 26086
rect 23484 25050 23540 25052
rect 23564 25050 23620 25052
rect 23644 25050 23700 25052
rect 23724 25050 23780 25052
rect 23484 24998 23530 25050
rect 23530 24998 23540 25050
rect 23564 24998 23594 25050
rect 23594 24998 23606 25050
rect 23606 24998 23620 25050
rect 23644 24998 23658 25050
rect 23658 24998 23670 25050
rect 23670 24998 23700 25050
rect 23724 24998 23734 25050
rect 23734 24998 23780 25050
rect 23484 24996 23540 24998
rect 23564 24996 23620 24998
rect 23644 24996 23700 24998
rect 23724 24996 23780 24998
rect 23484 23962 23540 23964
rect 23564 23962 23620 23964
rect 23644 23962 23700 23964
rect 23724 23962 23780 23964
rect 23484 23910 23530 23962
rect 23530 23910 23540 23962
rect 23564 23910 23594 23962
rect 23594 23910 23606 23962
rect 23606 23910 23620 23962
rect 23644 23910 23658 23962
rect 23658 23910 23670 23962
rect 23670 23910 23700 23962
rect 23724 23910 23734 23962
rect 23734 23910 23780 23962
rect 23484 23908 23540 23910
rect 23564 23908 23620 23910
rect 23644 23908 23700 23910
rect 23724 23908 23780 23910
rect 23484 22874 23540 22876
rect 23564 22874 23620 22876
rect 23644 22874 23700 22876
rect 23724 22874 23780 22876
rect 23484 22822 23530 22874
rect 23530 22822 23540 22874
rect 23564 22822 23594 22874
rect 23594 22822 23606 22874
rect 23606 22822 23620 22874
rect 23644 22822 23658 22874
rect 23658 22822 23670 22874
rect 23670 22822 23700 22874
rect 23724 22822 23734 22874
rect 23734 22822 23780 22874
rect 23484 22820 23540 22822
rect 23564 22820 23620 22822
rect 23644 22820 23700 22822
rect 23724 22820 23780 22822
rect 23484 21786 23540 21788
rect 23564 21786 23620 21788
rect 23644 21786 23700 21788
rect 23724 21786 23780 21788
rect 23484 21734 23530 21786
rect 23530 21734 23540 21786
rect 23564 21734 23594 21786
rect 23594 21734 23606 21786
rect 23606 21734 23620 21786
rect 23644 21734 23658 21786
rect 23658 21734 23670 21786
rect 23670 21734 23700 21786
rect 23724 21734 23734 21786
rect 23734 21734 23780 21786
rect 23484 21732 23540 21734
rect 23564 21732 23620 21734
rect 23644 21732 23700 21734
rect 23724 21732 23780 21734
rect 23484 20698 23540 20700
rect 23564 20698 23620 20700
rect 23644 20698 23700 20700
rect 23724 20698 23780 20700
rect 23484 20646 23530 20698
rect 23530 20646 23540 20698
rect 23564 20646 23594 20698
rect 23594 20646 23606 20698
rect 23606 20646 23620 20698
rect 23644 20646 23658 20698
rect 23658 20646 23670 20698
rect 23670 20646 23700 20698
rect 23724 20646 23734 20698
rect 23734 20646 23780 20698
rect 23484 20644 23540 20646
rect 23564 20644 23620 20646
rect 23644 20644 23700 20646
rect 23724 20644 23780 20646
rect 23484 19610 23540 19612
rect 23564 19610 23620 19612
rect 23644 19610 23700 19612
rect 23724 19610 23780 19612
rect 23484 19558 23530 19610
rect 23530 19558 23540 19610
rect 23564 19558 23594 19610
rect 23594 19558 23606 19610
rect 23606 19558 23620 19610
rect 23644 19558 23658 19610
rect 23658 19558 23670 19610
rect 23670 19558 23700 19610
rect 23724 19558 23734 19610
rect 23734 19558 23780 19610
rect 23484 19556 23540 19558
rect 23564 19556 23620 19558
rect 23644 19556 23700 19558
rect 23724 19556 23780 19558
rect 23484 18522 23540 18524
rect 23564 18522 23620 18524
rect 23644 18522 23700 18524
rect 23724 18522 23780 18524
rect 23484 18470 23530 18522
rect 23530 18470 23540 18522
rect 23564 18470 23594 18522
rect 23594 18470 23606 18522
rect 23606 18470 23620 18522
rect 23644 18470 23658 18522
rect 23658 18470 23670 18522
rect 23670 18470 23700 18522
rect 23724 18470 23734 18522
rect 23734 18470 23780 18522
rect 23484 18468 23540 18470
rect 23564 18468 23620 18470
rect 23644 18468 23700 18470
rect 23724 18468 23780 18470
rect 23484 17434 23540 17436
rect 23564 17434 23620 17436
rect 23644 17434 23700 17436
rect 23724 17434 23780 17436
rect 23484 17382 23530 17434
rect 23530 17382 23540 17434
rect 23564 17382 23594 17434
rect 23594 17382 23606 17434
rect 23606 17382 23620 17434
rect 23644 17382 23658 17434
rect 23658 17382 23670 17434
rect 23670 17382 23700 17434
rect 23724 17382 23734 17434
rect 23734 17382 23780 17434
rect 23484 17380 23540 17382
rect 23564 17380 23620 17382
rect 23644 17380 23700 17382
rect 23724 17380 23780 17382
rect 23484 16346 23540 16348
rect 23564 16346 23620 16348
rect 23644 16346 23700 16348
rect 23724 16346 23780 16348
rect 23484 16294 23530 16346
rect 23530 16294 23540 16346
rect 23564 16294 23594 16346
rect 23594 16294 23606 16346
rect 23606 16294 23620 16346
rect 23644 16294 23658 16346
rect 23658 16294 23670 16346
rect 23670 16294 23700 16346
rect 23724 16294 23734 16346
rect 23734 16294 23780 16346
rect 23484 16292 23540 16294
rect 23564 16292 23620 16294
rect 23644 16292 23700 16294
rect 23724 16292 23780 16294
rect 23484 15258 23540 15260
rect 23564 15258 23620 15260
rect 23644 15258 23700 15260
rect 23724 15258 23780 15260
rect 23484 15206 23530 15258
rect 23530 15206 23540 15258
rect 23564 15206 23594 15258
rect 23594 15206 23606 15258
rect 23606 15206 23620 15258
rect 23644 15206 23658 15258
rect 23658 15206 23670 15258
rect 23670 15206 23700 15258
rect 23724 15206 23734 15258
rect 23734 15206 23780 15258
rect 23484 15204 23540 15206
rect 23564 15204 23620 15206
rect 23644 15204 23700 15206
rect 23724 15204 23780 15206
rect 23484 14170 23540 14172
rect 23564 14170 23620 14172
rect 23644 14170 23700 14172
rect 23724 14170 23780 14172
rect 23484 14118 23530 14170
rect 23530 14118 23540 14170
rect 23564 14118 23594 14170
rect 23594 14118 23606 14170
rect 23606 14118 23620 14170
rect 23644 14118 23658 14170
rect 23658 14118 23670 14170
rect 23670 14118 23700 14170
rect 23724 14118 23734 14170
rect 23734 14118 23780 14170
rect 23484 14116 23540 14118
rect 23564 14116 23620 14118
rect 23644 14116 23700 14118
rect 23724 14116 23780 14118
rect 23484 13082 23540 13084
rect 23564 13082 23620 13084
rect 23644 13082 23700 13084
rect 23724 13082 23780 13084
rect 23484 13030 23530 13082
rect 23530 13030 23540 13082
rect 23564 13030 23594 13082
rect 23594 13030 23606 13082
rect 23606 13030 23620 13082
rect 23644 13030 23658 13082
rect 23658 13030 23670 13082
rect 23670 13030 23700 13082
rect 23724 13030 23734 13082
rect 23734 13030 23780 13082
rect 23484 13028 23540 13030
rect 23564 13028 23620 13030
rect 23644 13028 23700 13030
rect 23724 13028 23780 13030
rect 23484 11994 23540 11996
rect 23564 11994 23620 11996
rect 23644 11994 23700 11996
rect 23724 11994 23780 11996
rect 23484 11942 23530 11994
rect 23530 11942 23540 11994
rect 23564 11942 23594 11994
rect 23594 11942 23606 11994
rect 23606 11942 23620 11994
rect 23644 11942 23658 11994
rect 23658 11942 23670 11994
rect 23670 11942 23700 11994
rect 23724 11942 23734 11994
rect 23734 11942 23780 11994
rect 23484 11940 23540 11942
rect 23564 11940 23620 11942
rect 23644 11940 23700 11942
rect 23724 11940 23780 11942
rect 23484 10906 23540 10908
rect 23564 10906 23620 10908
rect 23644 10906 23700 10908
rect 23724 10906 23780 10908
rect 23484 10854 23530 10906
rect 23530 10854 23540 10906
rect 23564 10854 23594 10906
rect 23594 10854 23606 10906
rect 23606 10854 23620 10906
rect 23644 10854 23658 10906
rect 23658 10854 23670 10906
rect 23670 10854 23700 10906
rect 23724 10854 23734 10906
rect 23734 10854 23780 10906
rect 23484 10852 23540 10854
rect 23564 10852 23620 10854
rect 23644 10852 23700 10854
rect 23724 10852 23780 10854
rect 23484 9818 23540 9820
rect 23564 9818 23620 9820
rect 23644 9818 23700 9820
rect 23724 9818 23780 9820
rect 23484 9766 23530 9818
rect 23530 9766 23540 9818
rect 23564 9766 23594 9818
rect 23594 9766 23606 9818
rect 23606 9766 23620 9818
rect 23644 9766 23658 9818
rect 23658 9766 23670 9818
rect 23670 9766 23700 9818
rect 23724 9766 23734 9818
rect 23734 9766 23780 9818
rect 23484 9764 23540 9766
rect 23564 9764 23620 9766
rect 23644 9764 23700 9766
rect 23724 9764 23780 9766
rect 23484 8730 23540 8732
rect 23564 8730 23620 8732
rect 23644 8730 23700 8732
rect 23724 8730 23780 8732
rect 23484 8678 23530 8730
rect 23530 8678 23540 8730
rect 23564 8678 23594 8730
rect 23594 8678 23606 8730
rect 23606 8678 23620 8730
rect 23644 8678 23658 8730
rect 23658 8678 23670 8730
rect 23670 8678 23700 8730
rect 23724 8678 23734 8730
rect 23734 8678 23780 8730
rect 23484 8676 23540 8678
rect 23564 8676 23620 8678
rect 23644 8676 23700 8678
rect 23724 8676 23780 8678
rect 23484 7642 23540 7644
rect 23564 7642 23620 7644
rect 23644 7642 23700 7644
rect 23724 7642 23780 7644
rect 23484 7590 23530 7642
rect 23530 7590 23540 7642
rect 23564 7590 23594 7642
rect 23594 7590 23606 7642
rect 23606 7590 23620 7642
rect 23644 7590 23658 7642
rect 23658 7590 23670 7642
rect 23670 7590 23700 7642
rect 23724 7590 23734 7642
rect 23734 7590 23780 7642
rect 23484 7588 23540 7590
rect 23564 7588 23620 7590
rect 23644 7588 23700 7590
rect 23724 7588 23780 7590
rect 23484 6554 23540 6556
rect 23564 6554 23620 6556
rect 23644 6554 23700 6556
rect 23724 6554 23780 6556
rect 23484 6502 23530 6554
rect 23530 6502 23540 6554
rect 23564 6502 23594 6554
rect 23594 6502 23606 6554
rect 23606 6502 23620 6554
rect 23644 6502 23658 6554
rect 23658 6502 23670 6554
rect 23670 6502 23700 6554
rect 23724 6502 23734 6554
rect 23734 6502 23780 6554
rect 23484 6500 23540 6502
rect 23564 6500 23620 6502
rect 23644 6500 23700 6502
rect 23724 6500 23780 6502
rect 23484 5466 23540 5468
rect 23564 5466 23620 5468
rect 23644 5466 23700 5468
rect 23724 5466 23780 5468
rect 23484 5414 23530 5466
rect 23530 5414 23540 5466
rect 23564 5414 23594 5466
rect 23594 5414 23606 5466
rect 23606 5414 23620 5466
rect 23644 5414 23658 5466
rect 23658 5414 23670 5466
rect 23670 5414 23700 5466
rect 23724 5414 23734 5466
rect 23734 5414 23780 5466
rect 23484 5412 23540 5414
rect 23564 5412 23620 5414
rect 23644 5412 23700 5414
rect 23724 5412 23780 5414
rect 23484 4378 23540 4380
rect 23564 4378 23620 4380
rect 23644 4378 23700 4380
rect 23724 4378 23780 4380
rect 23484 4326 23530 4378
rect 23530 4326 23540 4378
rect 23564 4326 23594 4378
rect 23594 4326 23606 4378
rect 23606 4326 23620 4378
rect 23644 4326 23658 4378
rect 23658 4326 23670 4378
rect 23670 4326 23700 4378
rect 23724 4326 23734 4378
rect 23734 4326 23780 4378
rect 23484 4324 23540 4326
rect 23564 4324 23620 4326
rect 23644 4324 23700 4326
rect 23724 4324 23780 4326
rect 23484 3290 23540 3292
rect 23564 3290 23620 3292
rect 23644 3290 23700 3292
rect 23724 3290 23780 3292
rect 23484 3238 23530 3290
rect 23530 3238 23540 3290
rect 23564 3238 23594 3290
rect 23594 3238 23606 3290
rect 23606 3238 23620 3290
rect 23644 3238 23658 3290
rect 23658 3238 23670 3290
rect 23670 3238 23700 3290
rect 23724 3238 23734 3290
rect 23734 3238 23780 3290
rect 23484 3236 23540 3238
rect 23564 3236 23620 3238
rect 23644 3236 23700 3238
rect 23724 3236 23780 3238
rect 23484 2202 23540 2204
rect 23564 2202 23620 2204
rect 23644 2202 23700 2204
rect 23724 2202 23780 2204
rect 23484 2150 23530 2202
rect 23530 2150 23540 2202
rect 23564 2150 23594 2202
rect 23594 2150 23606 2202
rect 23606 2150 23620 2202
rect 23644 2150 23658 2202
rect 23658 2150 23670 2202
rect 23670 2150 23700 2202
rect 23724 2150 23734 2202
rect 23734 2150 23780 2202
rect 23484 2148 23540 2150
rect 23564 2148 23620 2150
rect 23644 2148 23700 2150
rect 23724 2148 23780 2150
rect 29116 33210 29172 33212
rect 29196 33210 29252 33212
rect 29276 33210 29332 33212
rect 29356 33210 29412 33212
rect 29116 33158 29162 33210
rect 29162 33158 29172 33210
rect 29196 33158 29226 33210
rect 29226 33158 29238 33210
rect 29238 33158 29252 33210
rect 29276 33158 29290 33210
rect 29290 33158 29302 33210
rect 29302 33158 29332 33210
rect 29356 33158 29366 33210
rect 29366 33158 29412 33210
rect 29116 33156 29172 33158
rect 29196 33156 29252 33158
rect 29276 33156 29332 33158
rect 29356 33156 29412 33158
rect 29116 32122 29172 32124
rect 29196 32122 29252 32124
rect 29276 32122 29332 32124
rect 29356 32122 29412 32124
rect 29116 32070 29162 32122
rect 29162 32070 29172 32122
rect 29196 32070 29226 32122
rect 29226 32070 29238 32122
rect 29238 32070 29252 32122
rect 29276 32070 29290 32122
rect 29290 32070 29302 32122
rect 29302 32070 29332 32122
rect 29356 32070 29366 32122
rect 29366 32070 29412 32122
rect 29116 32068 29172 32070
rect 29196 32068 29252 32070
rect 29276 32068 29332 32070
rect 29356 32068 29412 32070
rect 29116 31034 29172 31036
rect 29196 31034 29252 31036
rect 29276 31034 29332 31036
rect 29356 31034 29412 31036
rect 29116 30982 29162 31034
rect 29162 30982 29172 31034
rect 29196 30982 29226 31034
rect 29226 30982 29238 31034
rect 29238 30982 29252 31034
rect 29276 30982 29290 31034
rect 29290 30982 29302 31034
rect 29302 30982 29332 31034
rect 29356 30982 29366 31034
rect 29366 30982 29412 31034
rect 29116 30980 29172 30982
rect 29196 30980 29252 30982
rect 29276 30980 29332 30982
rect 29356 30980 29412 30982
rect 29116 29946 29172 29948
rect 29196 29946 29252 29948
rect 29276 29946 29332 29948
rect 29356 29946 29412 29948
rect 29116 29894 29162 29946
rect 29162 29894 29172 29946
rect 29196 29894 29226 29946
rect 29226 29894 29238 29946
rect 29238 29894 29252 29946
rect 29276 29894 29290 29946
rect 29290 29894 29302 29946
rect 29302 29894 29332 29946
rect 29356 29894 29366 29946
rect 29366 29894 29412 29946
rect 29116 29892 29172 29894
rect 29196 29892 29252 29894
rect 29276 29892 29332 29894
rect 29356 29892 29412 29894
rect 29116 28858 29172 28860
rect 29196 28858 29252 28860
rect 29276 28858 29332 28860
rect 29356 28858 29412 28860
rect 29116 28806 29162 28858
rect 29162 28806 29172 28858
rect 29196 28806 29226 28858
rect 29226 28806 29238 28858
rect 29238 28806 29252 28858
rect 29276 28806 29290 28858
rect 29290 28806 29302 28858
rect 29302 28806 29332 28858
rect 29356 28806 29366 28858
rect 29366 28806 29412 28858
rect 29116 28804 29172 28806
rect 29196 28804 29252 28806
rect 29276 28804 29332 28806
rect 29356 28804 29412 28806
rect 29116 27770 29172 27772
rect 29196 27770 29252 27772
rect 29276 27770 29332 27772
rect 29356 27770 29412 27772
rect 29116 27718 29162 27770
rect 29162 27718 29172 27770
rect 29196 27718 29226 27770
rect 29226 27718 29238 27770
rect 29238 27718 29252 27770
rect 29276 27718 29290 27770
rect 29290 27718 29302 27770
rect 29302 27718 29332 27770
rect 29356 27718 29366 27770
rect 29366 27718 29412 27770
rect 29116 27716 29172 27718
rect 29196 27716 29252 27718
rect 29276 27716 29332 27718
rect 29356 27716 29412 27718
rect 29116 26682 29172 26684
rect 29196 26682 29252 26684
rect 29276 26682 29332 26684
rect 29356 26682 29412 26684
rect 29116 26630 29162 26682
rect 29162 26630 29172 26682
rect 29196 26630 29226 26682
rect 29226 26630 29238 26682
rect 29238 26630 29252 26682
rect 29276 26630 29290 26682
rect 29290 26630 29302 26682
rect 29302 26630 29332 26682
rect 29356 26630 29366 26682
rect 29366 26630 29412 26682
rect 29116 26628 29172 26630
rect 29196 26628 29252 26630
rect 29276 26628 29332 26630
rect 29356 26628 29412 26630
rect 29116 25594 29172 25596
rect 29196 25594 29252 25596
rect 29276 25594 29332 25596
rect 29356 25594 29412 25596
rect 29116 25542 29162 25594
rect 29162 25542 29172 25594
rect 29196 25542 29226 25594
rect 29226 25542 29238 25594
rect 29238 25542 29252 25594
rect 29276 25542 29290 25594
rect 29290 25542 29302 25594
rect 29302 25542 29332 25594
rect 29356 25542 29366 25594
rect 29366 25542 29412 25594
rect 29116 25540 29172 25542
rect 29196 25540 29252 25542
rect 29276 25540 29332 25542
rect 29356 25540 29412 25542
rect 29116 24506 29172 24508
rect 29196 24506 29252 24508
rect 29276 24506 29332 24508
rect 29356 24506 29412 24508
rect 29116 24454 29162 24506
rect 29162 24454 29172 24506
rect 29196 24454 29226 24506
rect 29226 24454 29238 24506
rect 29238 24454 29252 24506
rect 29276 24454 29290 24506
rect 29290 24454 29302 24506
rect 29302 24454 29332 24506
rect 29356 24454 29366 24506
rect 29366 24454 29412 24506
rect 29116 24452 29172 24454
rect 29196 24452 29252 24454
rect 29276 24452 29332 24454
rect 29356 24452 29412 24454
rect 29116 23418 29172 23420
rect 29196 23418 29252 23420
rect 29276 23418 29332 23420
rect 29356 23418 29412 23420
rect 29116 23366 29162 23418
rect 29162 23366 29172 23418
rect 29196 23366 29226 23418
rect 29226 23366 29238 23418
rect 29238 23366 29252 23418
rect 29276 23366 29290 23418
rect 29290 23366 29302 23418
rect 29302 23366 29332 23418
rect 29356 23366 29366 23418
rect 29366 23366 29412 23418
rect 29116 23364 29172 23366
rect 29196 23364 29252 23366
rect 29276 23364 29332 23366
rect 29356 23364 29412 23366
rect 29116 22330 29172 22332
rect 29196 22330 29252 22332
rect 29276 22330 29332 22332
rect 29356 22330 29412 22332
rect 29116 22278 29162 22330
rect 29162 22278 29172 22330
rect 29196 22278 29226 22330
rect 29226 22278 29238 22330
rect 29238 22278 29252 22330
rect 29276 22278 29290 22330
rect 29290 22278 29302 22330
rect 29302 22278 29332 22330
rect 29356 22278 29366 22330
rect 29366 22278 29412 22330
rect 29116 22276 29172 22278
rect 29196 22276 29252 22278
rect 29276 22276 29332 22278
rect 29356 22276 29412 22278
rect 29116 21242 29172 21244
rect 29196 21242 29252 21244
rect 29276 21242 29332 21244
rect 29356 21242 29412 21244
rect 29116 21190 29162 21242
rect 29162 21190 29172 21242
rect 29196 21190 29226 21242
rect 29226 21190 29238 21242
rect 29238 21190 29252 21242
rect 29276 21190 29290 21242
rect 29290 21190 29302 21242
rect 29302 21190 29332 21242
rect 29356 21190 29366 21242
rect 29366 21190 29412 21242
rect 29116 21188 29172 21190
rect 29196 21188 29252 21190
rect 29276 21188 29332 21190
rect 29356 21188 29412 21190
rect 29116 20154 29172 20156
rect 29196 20154 29252 20156
rect 29276 20154 29332 20156
rect 29356 20154 29412 20156
rect 29116 20102 29162 20154
rect 29162 20102 29172 20154
rect 29196 20102 29226 20154
rect 29226 20102 29238 20154
rect 29238 20102 29252 20154
rect 29276 20102 29290 20154
rect 29290 20102 29302 20154
rect 29302 20102 29332 20154
rect 29356 20102 29366 20154
rect 29366 20102 29412 20154
rect 29116 20100 29172 20102
rect 29196 20100 29252 20102
rect 29276 20100 29332 20102
rect 29356 20100 29412 20102
rect 29116 19066 29172 19068
rect 29196 19066 29252 19068
rect 29276 19066 29332 19068
rect 29356 19066 29412 19068
rect 29116 19014 29162 19066
rect 29162 19014 29172 19066
rect 29196 19014 29226 19066
rect 29226 19014 29238 19066
rect 29238 19014 29252 19066
rect 29276 19014 29290 19066
rect 29290 19014 29302 19066
rect 29302 19014 29332 19066
rect 29356 19014 29366 19066
rect 29366 19014 29412 19066
rect 29116 19012 29172 19014
rect 29196 19012 29252 19014
rect 29276 19012 29332 19014
rect 29356 19012 29412 19014
rect 29116 17978 29172 17980
rect 29196 17978 29252 17980
rect 29276 17978 29332 17980
rect 29356 17978 29412 17980
rect 29116 17926 29162 17978
rect 29162 17926 29172 17978
rect 29196 17926 29226 17978
rect 29226 17926 29238 17978
rect 29238 17926 29252 17978
rect 29276 17926 29290 17978
rect 29290 17926 29302 17978
rect 29302 17926 29332 17978
rect 29356 17926 29366 17978
rect 29366 17926 29412 17978
rect 29116 17924 29172 17926
rect 29196 17924 29252 17926
rect 29276 17924 29332 17926
rect 29356 17924 29412 17926
rect 33138 33360 33194 33416
rect 33782 35400 33838 35456
rect 33690 34040 33746 34096
rect 34242 34720 34298 34776
rect 34242 32000 34298 32056
rect 29116 16890 29172 16892
rect 29196 16890 29252 16892
rect 29276 16890 29332 16892
rect 29356 16890 29412 16892
rect 29116 16838 29162 16890
rect 29162 16838 29172 16890
rect 29196 16838 29226 16890
rect 29226 16838 29238 16890
rect 29238 16838 29252 16890
rect 29276 16838 29290 16890
rect 29290 16838 29302 16890
rect 29302 16838 29332 16890
rect 29356 16838 29366 16890
rect 29366 16838 29412 16890
rect 29116 16836 29172 16838
rect 29196 16836 29252 16838
rect 29276 16836 29332 16838
rect 29356 16836 29412 16838
rect 29116 15802 29172 15804
rect 29196 15802 29252 15804
rect 29276 15802 29332 15804
rect 29356 15802 29412 15804
rect 29116 15750 29162 15802
rect 29162 15750 29172 15802
rect 29196 15750 29226 15802
rect 29226 15750 29238 15802
rect 29238 15750 29252 15802
rect 29276 15750 29290 15802
rect 29290 15750 29302 15802
rect 29302 15750 29332 15802
rect 29356 15750 29366 15802
rect 29366 15750 29412 15802
rect 29116 15748 29172 15750
rect 29196 15748 29252 15750
rect 29276 15748 29332 15750
rect 29356 15748 29412 15750
rect 29116 14714 29172 14716
rect 29196 14714 29252 14716
rect 29276 14714 29332 14716
rect 29356 14714 29412 14716
rect 29116 14662 29162 14714
rect 29162 14662 29172 14714
rect 29196 14662 29226 14714
rect 29226 14662 29238 14714
rect 29238 14662 29252 14714
rect 29276 14662 29290 14714
rect 29290 14662 29302 14714
rect 29302 14662 29332 14714
rect 29356 14662 29366 14714
rect 29366 14662 29412 14714
rect 29116 14660 29172 14662
rect 29196 14660 29252 14662
rect 29276 14660 29332 14662
rect 29356 14660 29412 14662
rect 29116 13626 29172 13628
rect 29196 13626 29252 13628
rect 29276 13626 29332 13628
rect 29356 13626 29412 13628
rect 29116 13574 29162 13626
rect 29162 13574 29172 13626
rect 29196 13574 29226 13626
rect 29226 13574 29238 13626
rect 29238 13574 29252 13626
rect 29276 13574 29290 13626
rect 29290 13574 29302 13626
rect 29302 13574 29332 13626
rect 29356 13574 29366 13626
rect 29366 13574 29412 13626
rect 29116 13572 29172 13574
rect 29196 13572 29252 13574
rect 29276 13572 29332 13574
rect 29356 13572 29412 13574
rect 29116 12538 29172 12540
rect 29196 12538 29252 12540
rect 29276 12538 29332 12540
rect 29356 12538 29412 12540
rect 29116 12486 29162 12538
rect 29162 12486 29172 12538
rect 29196 12486 29226 12538
rect 29226 12486 29238 12538
rect 29238 12486 29252 12538
rect 29276 12486 29290 12538
rect 29290 12486 29302 12538
rect 29302 12486 29332 12538
rect 29356 12486 29366 12538
rect 29366 12486 29412 12538
rect 29116 12484 29172 12486
rect 29196 12484 29252 12486
rect 29276 12484 29332 12486
rect 29356 12484 29412 12486
rect 29116 11450 29172 11452
rect 29196 11450 29252 11452
rect 29276 11450 29332 11452
rect 29356 11450 29412 11452
rect 29116 11398 29162 11450
rect 29162 11398 29172 11450
rect 29196 11398 29226 11450
rect 29226 11398 29238 11450
rect 29238 11398 29252 11450
rect 29276 11398 29290 11450
rect 29290 11398 29302 11450
rect 29302 11398 29332 11450
rect 29356 11398 29366 11450
rect 29366 11398 29412 11450
rect 29116 11396 29172 11398
rect 29196 11396 29252 11398
rect 29276 11396 29332 11398
rect 29356 11396 29412 11398
rect 29116 10362 29172 10364
rect 29196 10362 29252 10364
rect 29276 10362 29332 10364
rect 29356 10362 29412 10364
rect 29116 10310 29162 10362
rect 29162 10310 29172 10362
rect 29196 10310 29226 10362
rect 29226 10310 29238 10362
rect 29238 10310 29252 10362
rect 29276 10310 29290 10362
rect 29290 10310 29302 10362
rect 29302 10310 29332 10362
rect 29356 10310 29366 10362
rect 29366 10310 29412 10362
rect 29116 10308 29172 10310
rect 29196 10308 29252 10310
rect 29276 10308 29332 10310
rect 29356 10308 29412 10310
rect 29116 9274 29172 9276
rect 29196 9274 29252 9276
rect 29276 9274 29332 9276
rect 29356 9274 29412 9276
rect 29116 9222 29162 9274
rect 29162 9222 29172 9274
rect 29196 9222 29226 9274
rect 29226 9222 29238 9274
rect 29238 9222 29252 9274
rect 29276 9222 29290 9274
rect 29290 9222 29302 9274
rect 29302 9222 29332 9274
rect 29356 9222 29366 9274
rect 29366 9222 29412 9274
rect 29116 9220 29172 9222
rect 29196 9220 29252 9222
rect 29276 9220 29332 9222
rect 29356 9220 29412 9222
rect 29116 8186 29172 8188
rect 29196 8186 29252 8188
rect 29276 8186 29332 8188
rect 29356 8186 29412 8188
rect 29116 8134 29162 8186
rect 29162 8134 29172 8186
rect 29196 8134 29226 8186
rect 29226 8134 29238 8186
rect 29238 8134 29252 8186
rect 29276 8134 29290 8186
rect 29290 8134 29302 8186
rect 29302 8134 29332 8186
rect 29356 8134 29366 8186
rect 29366 8134 29412 8186
rect 29116 8132 29172 8134
rect 29196 8132 29252 8134
rect 29276 8132 29332 8134
rect 29356 8132 29412 8134
rect 29116 7098 29172 7100
rect 29196 7098 29252 7100
rect 29276 7098 29332 7100
rect 29356 7098 29412 7100
rect 29116 7046 29162 7098
rect 29162 7046 29172 7098
rect 29196 7046 29226 7098
rect 29226 7046 29238 7098
rect 29238 7046 29252 7098
rect 29276 7046 29290 7098
rect 29290 7046 29302 7098
rect 29302 7046 29332 7098
rect 29356 7046 29366 7098
rect 29366 7046 29412 7098
rect 29116 7044 29172 7046
rect 29196 7044 29252 7046
rect 29276 7044 29332 7046
rect 29356 7044 29412 7046
rect 29116 6010 29172 6012
rect 29196 6010 29252 6012
rect 29276 6010 29332 6012
rect 29356 6010 29412 6012
rect 29116 5958 29162 6010
rect 29162 5958 29172 6010
rect 29196 5958 29226 6010
rect 29226 5958 29238 6010
rect 29238 5958 29252 6010
rect 29276 5958 29290 6010
rect 29290 5958 29302 6010
rect 29302 5958 29332 6010
rect 29356 5958 29366 6010
rect 29366 5958 29412 6010
rect 29116 5956 29172 5958
rect 29196 5956 29252 5958
rect 29276 5956 29332 5958
rect 29356 5956 29412 5958
rect 29116 4922 29172 4924
rect 29196 4922 29252 4924
rect 29276 4922 29332 4924
rect 29356 4922 29412 4924
rect 29116 4870 29162 4922
rect 29162 4870 29172 4922
rect 29196 4870 29226 4922
rect 29226 4870 29238 4922
rect 29238 4870 29252 4922
rect 29276 4870 29290 4922
rect 29290 4870 29302 4922
rect 29302 4870 29332 4922
rect 29356 4870 29366 4922
rect 29366 4870 29412 4922
rect 29116 4868 29172 4870
rect 29196 4868 29252 4870
rect 29276 4868 29332 4870
rect 29356 4868 29412 4870
rect 29116 3834 29172 3836
rect 29196 3834 29252 3836
rect 29276 3834 29332 3836
rect 29356 3834 29412 3836
rect 29116 3782 29162 3834
rect 29162 3782 29172 3834
rect 29196 3782 29226 3834
rect 29226 3782 29238 3834
rect 29238 3782 29252 3834
rect 29276 3782 29290 3834
rect 29290 3782 29302 3834
rect 29302 3782 29332 3834
rect 29356 3782 29366 3834
rect 29366 3782 29412 3834
rect 29116 3780 29172 3782
rect 29196 3780 29252 3782
rect 29276 3780 29332 3782
rect 29356 3780 29412 3782
rect 29116 2746 29172 2748
rect 29196 2746 29252 2748
rect 29276 2746 29332 2748
rect 29356 2746 29412 2748
rect 29116 2694 29162 2746
rect 29162 2694 29172 2746
rect 29196 2694 29226 2746
rect 29226 2694 29238 2746
rect 29238 2694 29252 2746
rect 29276 2694 29290 2746
rect 29290 2694 29302 2746
rect 29302 2694 29332 2746
rect 29356 2694 29366 2746
rect 29366 2694 29412 2746
rect 29116 2692 29172 2694
rect 29196 2692 29252 2694
rect 29276 2692 29332 2694
rect 29356 2692 29412 2694
rect 34334 31340 34390 31376
rect 34334 31320 34336 31340
rect 34336 31320 34388 31340
rect 34388 31320 34390 31340
rect 33506 20440 33562 20496
rect 34334 30676 34336 30696
rect 34336 30676 34388 30696
rect 34388 30676 34390 30696
rect 34334 30640 34390 30676
rect 34334 29960 34390 30016
rect 34334 29280 34390 29336
rect 34242 28600 34298 28656
rect 34242 27940 34298 27976
rect 34242 27920 34244 27940
rect 34244 27920 34296 27940
rect 34296 27920 34298 27940
rect 32402 3476 32404 3496
rect 32404 3476 32456 3496
rect 32456 3476 32458 3496
rect 32402 3440 32458 3476
rect 32586 2080 32642 2136
rect 34242 26560 34298 26616
rect 34334 25880 34390 25936
rect 34242 25200 34298 25256
rect 34242 24556 34244 24576
rect 34244 24556 34296 24576
rect 34296 24556 34298 24576
rect 34242 24520 34298 24556
rect 34242 23840 34298 23896
rect 34242 23196 34244 23216
rect 34244 23196 34296 23216
rect 34296 23196 34298 23216
rect 34242 23160 34298 23196
rect 34334 22516 34336 22536
rect 34336 22516 34388 22536
rect 34388 22516 34390 22536
rect 34334 22480 34390 22516
rect 34334 21120 34390 21176
rect 34334 19796 34336 19816
rect 34336 19796 34388 19816
rect 34388 19796 34390 19816
rect 34334 19760 34390 19796
rect 34334 19080 34390 19136
rect 34334 18400 34390 18456
rect 34242 17720 34298 17776
rect 34242 17060 34298 17096
rect 34242 17040 34244 17060
rect 34244 17040 34296 17060
rect 34296 17040 34298 17060
rect 34334 15680 34390 15736
rect 34242 15000 34298 15056
rect 34334 14356 34336 14376
rect 34336 14356 34388 14376
rect 34388 14356 34390 14376
rect 34334 14320 34390 14356
rect 34334 13640 34390 13696
rect 34242 12960 34298 13016
rect 34242 12280 34298 12336
rect 34242 11620 34298 11656
rect 34242 11600 34244 11620
rect 34244 11600 34296 11620
rect 34296 11600 34298 11620
rect 34334 9560 34390 9616
rect 34242 8880 34298 8936
rect 34242 8200 34298 8256
rect 34242 7520 34298 7576
rect 34242 6840 34298 6896
rect 34242 6160 34298 6216
rect 34334 4800 34390 4856
rect 34242 4120 34298 4176
rect 33138 1400 33194 1456
rect 34242 2760 34298 2816
rect 33874 720 33930 776
<< metal3 >>
rect 0 35458 800 35488
rect 2957 35458 3023 35461
rect 0 35456 3023 35458
rect 0 35400 2962 35456
rect 3018 35400 3023 35456
rect 0 35398 3023 35400
rect 0 35368 800 35398
rect 2957 35395 3023 35398
rect 33777 35458 33843 35461
rect 35200 35458 36000 35488
rect 33777 35456 36000 35458
rect 33777 35400 33782 35456
rect 33838 35400 36000 35456
rect 33777 35398 36000 35400
rect 33777 35395 33843 35398
rect 35200 35368 36000 35398
rect 0 34778 800 34808
rect 2865 34778 2931 34781
rect 0 34776 2931 34778
rect 0 34720 2870 34776
rect 2926 34720 2931 34776
rect 0 34718 2931 34720
rect 0 34688 800 34718
rect 2865 34715 2931 34718
rect 34237 34778 34303 34781
rect 35200 34778 36000 34808
rect 34237 34776 36000 34778
rect 34237 34720 34242 34776
rect 34298 34720 36000 34776
rect 34237 34718 36000 34720
rect 34237 34715 34303 34718
rect 35200 34688 36000 34718
rect 0 34098 800 34128
rect 2129 34098 2195 34101
rect 0 34096 2195 34098
rect 0 34040 2134 34096
rect 2190 34040 2195 34096
rect 0 34038 2195 34040
rect 0 34008 800 34038
rect 2129 34035 2195 34038
rect 33685 34098 33751 34101
rect 35200 34098 36000 34128
rect 33685 34096 36000 34098
rect 33685 34040 33690 34096
rect 33746 34040 36000 34096
rect 33685 34038 36000 34040
rect 33685 34035 33751 34038
rect 35200 34008 36000 34038
rect 12208 33760 12528 33761
rect 12208 33696 12216 33760
rect 12280 33696 12296 33760
rect 12360 33696 12376 33760
rect 12440 33696 12456 33760
rect 12520 33696 12528 33760
rect 12208 33695 12528 33696
rect 23472 33760 23792 33761
rect 23472 33696 23480 33760
rect 23544 33696 23560 33760
rect 23624 33696 23640 33760
rect 23704 33696 23720 33760
rect 23784 33696 23792 33760
rect 23472 33695 23792 33696
rect 0 33328 800 33448
rect 33133 33418 33199 33421
rect 35200 33418 36000 33448
rect 33133 33416 36000 33418
rect 33133 33360 33138 33416
rect 33194 33360 36000 33416
rect 33133 33358 36000 33360
rect 33133 33355 33199 33358
rect 35200 33328 36000 33358
rect 6576 33216 6896 33217
rect 6576 33152 6584 33216
rect 6648 33152 6664 33216
rect 6728 33152 6744 33216
rect 6808 33152 6824 33216
rect 6888 33152 6896 33216
rect 6576 33151 6896 33152
rect 17840 33216 18160 33217
rect 17840 33152 17848 33216
rect 17912 33152 17928 33216
rect 17992 33152 18008 33216
rect 18072 33152 18088 33216
rect 18152 33152 18160 33216
rect 17840 33151 18160 33152
rect 29104 33216 29424 33217
rect 29104 33152 29112 33216
rect 29176 33152 29192 33216
rect 29256 33152 29272 33216
rect 29336 33152 29352 33216
rect 29416 33152 29424 33216
rect 29104 33151 29424 33152
rect 12208 32672 12528 32673
rect 12208 32608 12216 32672
rect 12280 32608 12296 32672
rect 12360 32608 12376 32672
rect 12440 32608 12456 32672
rect 12520 32608 12528 32672
rect 12208 32607 12528 32608
rect 23472 32672 23792 32673
rect 23472 32608 23480 32672
rect 23544 32608 23560 32672
rect 23624 32608 23640 32672
rect 23704 32608 23720 32672
rect 23784 32608 23792 32672
rect 23472 32607 23792 32608
rect 6576 32128 6896 32129
rect 0 32058 800 32088
rect 6576 32064 6584 32128
rect 6648 32064 6664 32128
rect 6728 32064 6744 32128
rect 6808 32064 6824 32128
rect 6888 32064 6896 32128
rect 6576 32063 6896 32064
rect 17840 32128 18160 32129
rect 17840 32064 17848 32128
rect 17912 32064 17928 32128
rect 17992 32064 18008 32128
rect 18072 32064 18088 32128
rect 18152 32064 18160 32128
rect 17840 32063 18160 32064
rect 29104 32128 29424 32129
rect 29104 32064 29112 32128
rect 29176 32064 29192 32128
rect 29256 32064 29272 32128
rect 29336 32064 29352 32128
rect 29416 32064 29424 32128
rect 29104 32063 29424 32064
rect 1393 32058 1459 32061
rect 0 32056 1459 32058
rect 0 32000 1398 32056
rect 1454 32000 1459 32056
rect 0 31998 1459 32000
rect 0 31968 800 31998
rect 1393 31995 1459 31998
rect 34237 32058 34303 32061
rect 35200 32058 36000 32088
rect 34237 32056 36000 32058
rect 34237 32000 34242 32056
rect 34298 32000 36000 32056
rect 34237 31998 36000 32000
rect 34237 31995 34303 31998
rect 35200 31968 36000 31998
rect 1669 31922 1735 31925
rect 15285 31922 15351 31925
rect 1669 31920 15351 31922
rect 1669 31864 1674 31920
rect 1730 31864 15290 31920
rect 15346 31864 15351 31920
rect 1669 31862 15351 31864
rect 1669 31859 1735 31862
rect 15285 31859 15351 31862
rect 12208 31584 12528 31585
rect 12208 31520 12216 31584
rect 12280 31520 12296 31584
rect 12360 31520 12376 31584
rect 12440 31520 12456 31584
rect 12520 31520 12528 31584
rect 12208 31519 12528 31520
rect 23472 31584 23792 31585
rect 23472 31520 23480 31584
rect 23544 31520 23560 31584
rect 23624 31520 23640 31584
rect 23704 31520 23720 31584
rect 23784 31520 23792 31584
rect 23472 31519 23792 31520
rect 0 31378 800 31408
rect 1485 31378 1551 31381
rect 0 31376 1551 31378
rect 0 31320 1490 31376
rect 1546 31320 1551 31376
rect 0 31318 1551 31320
rect 0 31288 800 31318
rect 1485 31315 1551 31318
rect 34329 31378 34395 31381
rect 35200 31378 36000 31408
rect 34329 31376 36000 31378
rect 34329 31320 34334 31376
rect 34390 31320 36000 31376
rect 34329 31318 36000 31320
rect 34329 31315 34395 31318
rect 35200 31288 36000 31318
rect 6576 31040 6896 31041
rect 6576 30976 6584 31040
rect 6648 30976 6664 31040
rect 6728 30976 6744 31040
rect 6808 30976 6824 31040
rect 6888 30976 6896 31040
rect 6576 30975 6896 30976
rect 17840 31040 18160 31041
rect 17840 30976 17848 31040
rect 17912 30976 17928 31040
rect 17992 30976 18008 31040
rect 18072 30976 18088 31040
rect 18152 30976 18160 31040
rect 17840 30975 18160 30976
rect 29104 31040 29424 31041
rect 29104 30976 29112 31040
rect 29176 30976 29192 31040
rect 29256 30976 29272 31040
rect 29336 30976 29352 31040
rect 29416 30976 29424 31040
rect 29104 30975 29424 30976
rect 0 30698 800 30728
rect 1485 30698 1551 30701
rect 0 30696 1551 30698
rect 0 30640 1490 30696
rect 1546 30640 1551 30696
rect 0 30638 1551 30640
rect 0 30608 800 30638
rect 1485 30635 1551 30638
rect 34329 30698 34395 30701
rect 35200 30698 36000 30728
rect 34329 30696 36000 30698
rect 34329 30640 34334 30696
rect 34390 30640 36000 30696
rect 34329 30638 36000 30640
rect 34329 30635 34395 30638
rect 35200 30608 36000 30638
rect 12208 30496 12528 30497
rect 12208 30432 12216 30496
rect 12280 30432 12296 30496
rect 12360 30432 12376 30496
rect 12440 30432 12456 30496
rect 12520 30432 12528 30496
rect 12208 30431 12528 30432
rect 23472 30496 23792 30497
rect 23472 30432 23480 30496
rect 23544 30432 23560 30496
rect 23624 30432 23640 30496
rect 23704 30432 23720 30496
rect 23784 30432 23792 30496
rect 23472 30431 23792 30432
rect 0 30018 800 30048
rect 1945 30018 2011 30021
rect 0 30016 2011 30018
rect 0 29960 1950 30016
rect 2006 29960 2011 30016
rect 0 29958 2011 29960
rect 0 29928 800 29958
rect 1945 29955 2011 29958
rect 34329 30018 34395 30021
rect 35200 30018 36000 30048
rect 34329 30016 36000 30018
rect 34329 29960 34334 30016
rect 34390 29960 36000 30016
rect 34329 29958 36000 29960
rect 34329 29955 34395 29958
rect 6576 29952 6896 29953
rect 6576 29888 6584 29952
rect 6648 29888 6664 29952
rect 6728 29888 6744 29952
rect 6808 29888 6824 29952
rect 6888 29888 6896 29952
rect 6576 29887 6896 29888
rect 17840 29952 18160 29953
rect 17840 29888 17848 29952
rect 17912 29888 17928 29952
rect 17992 29888 18008 29952
rect 18072 29888 18088 29952
rect 18152 29888 18160 29952
rect 17840 29887 18160 29888
rect 29104 29952 29424 29953
rect 29104 29888 29112 29952
rect 29176 29888 29192 29952
rect 29256 29888 29272 29952
rect 29336 29888 29352 29952
rect 29416 29888 29424 29952
rect 35200 29928 36000 29958
rect 29104 29887 29424 29888
rect 12208 29408 12528 29409
rect 0 29338 800 29368
rect 12208 29344 12216 29408
rect 12280 29344 12296 29408
rect 12360 29344 12376 29408
rect 12440 29344 12456 29408
rect 12520 29344 12528 29408
rect 12208 29343 12528 29344
rect 23472 29408 23792 29409
rect 23472 29344 23480 29408
rect 23544 29344 23560 29408
rect 23624 29344 23640 29408
rect 23704 29344 23720 29408
rect 23784 29344 23792 29408
rect 23472 29343 23792 29344
rect 1485 29338 1551 29341
rect 0 29336 1551 29338
rect 0 29280 1490 29336
rect 1546 29280 1551 29336
rect 0 29278 1551 29280
rect 0 29248 800 29278
rect 1485 29275 1551 29278
rect 34329 29338 34395 29341
rect 35200 29338 36000 29368
rect 34329 29336 36000 29338
rect 34329 29280 34334 29336
rect 34390 29280 36000 29336
rect 34329 29278 36000 29280
rect 34329 29275 34395 29278
rect 35200 29248 36000 29278
rect 6576 28864 6896 28865
rect 6576 28800 6584 28864
rect 6648 28800 6664 28864
rect 6728 28800 6744 28864
rect 6808 28800 6824 28864
rect 6888 28800 6896 28864
rect 6576 28799 6896 28800
rect 17840 28864 18160 28865
rect 17840 28800 17848 28864
rect 17912 28800 17928 28864
rect 17992 28800 18008 28864
rect 18072 28800 18088 28864
rect 18152 28800 18160 28864
rect 17840 28799 18160 28800
rect 29104 28864 29424 28865
rect 29104 28800 29112 28864
rect 29176 28800 29192 28864
rect 29256 28800 29272 28864
rect 29336 28800 29352 28864
rect 29416 28800 29424 28864
rect 29104 28799 29424 28800
rect 0 28658 800 28688
rect 1669 28658 1735 28661
rect 0 28656 1735 28658
rect 0 28600 1674 28656
rect 1730 28600 1735 28656
rect 0 28598 1735 28600
rect 0 28568 800 28598
rect 1669 28595 1735 28598
rect 34237 28658 34303 28661
rect 35200 28658 36000 28688
rect 34237 28656 36000 28658
rect 34237 28600 34242 28656
rect 34298 28600 36000 28656
rect 34237 28598 36000 28600
rect 34237 28595 34303 28598
rect 35200 28568 36000 28598
rect 12208 28320 12528 28321
rect 12208 28256 12216 28320
rect 12280 28256 12296 28320
rect 12360 28256 12376 28320
rect 12440 28256 12456 28320
rect 12520 28256 12528 28320
rect 12208 28255 12528 28256
rect 23472 28320 23792 28321
rect 23472 28256 23480 28320
rect 23544 28256 23560 28320
rect 23624 28256 23640 28320
rect 23704 28256 23720 28320
rect 23784 28256 23792 28320
rect 23472 28255 23792 28256
rect 0 27978 800 28008
rect 1485 27978 1551 27981
rect 0 27976 1551 27978
rect 0 27920 1490 27976
rect 1546 27920 1551 27976
rect 0 27918 1551 27920
rect 0 27888 800 27918
rect 1485 27915 1551 27918
rect 34237 27978 34303 27981
rect 35200 27978 36000 28008
rect 34237 27976 36000 27978
rect 34237 27920 34242 27976
rect 34298 27920 36000 27976
rect 34237 27918 36000 27920
rect 34237 27915 34303 27918
rect 35200 27888 36000 27918
rect 6576 27776 6896 27777
rect 6576 27712 6584 27776
rect 6648 27712 6664 27776
rect 6728 27712 6744 27776
rect 6808 27712 6824 27776
rect 6888 27712 6896 27776
rect 6576 27711 6896 27712
rect 17840 27776 18160 27777
rect 17840 27712 17848 27776
rect 17912 27712 17928 27776
rect 17992 27712 18008 27776
rect 18072 27712 18088 27776
rect 18152 27712 18160 27776
rect 17840 27711 18160 27712
rect 29104 27776 29424 27777
rect 29104 27712 29112 27776
rect 29176 27712 29192 27776
rect 29256 27712 29272 27776
rect 29336 27712 29352 27776
rect 29416 27712 29424 27776
rect 29104 27711 29424 27712
rect 12208 27232 12528 27233
rect 12208 27168 12216 27232
rect 12280 27168 12296 27232
rect 12360 27168 12376 27232
rect 12440 27168 12456 27232
rect 12520 27168 12528 27232
rect 12208 27167 12528 27168
rect 23472 27232 23792 27233
rect 23472 27168 23480 27232
rect 23544 27168 23560 27232
rect 23624 27168 23640 27232
rect 23704 27168 23720 27232
rect 23784 27168 23792 27232
rect 23472 27167 23792 27168
rect 6576 26688 6896 26689
rect 0 26528 800 26648
rect 6576 26624 6584 26688
rect 6648 26624 6664 26688
rect 6728 26624 6744 26688
rect 6808 26624 6824 26688
rect 6888 26624 6896 26688
rect 6576 26623 6896 26624
rect 17840 26688 18160 26689
rect 17840 26624 17848 26688
rect 17912 26624 17928 26688
rect 17992 26624 18008 26688
rect 18072 26624 18088 26688
rect 18152 26624 18160 26688
rect 17840 26623 18160 26624
rect 29104 26688 29424 26689
rect 29104 26624 29112 26688
rect 29176 26624 29192 26688
rect 29256 26624 29272 26688
rect 29336 26624 29352 26688
rect 29416 26624 29424 26688
rect 29104 26623 29424 26624
rect 34237 26618 34303 26621
rect 35200 26618 36000 26648
rect 34237 26616 36000 26618
rect 34237 26560 34242 26616
rect 34298 26560 36000 26616
rect 34237 26558 36000 26560
rect 34237 26555 34303 26558
rect 35200 26528 36000 26558
rect 12208 26144 12528 26145
rect 12208 26080 12216 26144
rect 12280 26080 12296 26144
rect 12360 26080 12376 26144
rect 12440 26080 12456 26144
rect 12520 26080 12528 26144
rect 12208 26079 12528 26080
rect 23472 26144 23792 26145
rect 23472 26080 23480 26144
rect 23544 26080 23560 26144
rect 23624 26080 23640 26144
rect 23704 26080 23720 26144
rect 23784 26080 23792 26144
rect 23472 26079 23792 26080
rect 0 25938 800 25968
rect 1393 25938 1459 25941
rect 0 25936 1459 25938
rect 0 25880 1398 25936
rect 1454 25880 1459 25936
rect 0 25878 1459 25880
rect 0 25848 800 25878
rect 1393 25875 1459 25878
rect 34329 25938 34395 25941
rect 35200 25938 36000 25968
rect 34329 25936 36000 25938
rect 34329 25880 34334 25936
rect 34390 25880 36000 25936
rect 34329 25878 36000 25880
rect 34329 25875 34395 25878
rect 35200 25848 36000 25878
rect 6576 25600 6896 25601
rect 6576 25536 6584 25600
rect 6648 25536 6664 25600
rect 6728 25536 6744 25600
rect 6808 25536 6824 25600
rect 6888 25536 6896 25600
rect 6576 25535 6896 25536
rect 17840 25600 18160 25601
rect 17840 25536 17848 25600
rect 17912 25536 17928 25600
rect 17992 25536 18008 25600
rect 18072 25536 18088 25600
rect 18152 25536 18160 25600
rect 17840 25535 18160 25536
rect 29104 25600 29424 25601
rect 29104 25536 29112 25600
rect 29176 25536 29192 25600
rect 29256 25536 29272 25600
rect 29336 25536 29352 25600
rect 29416 25536 29424 25600
rect 29104 25535 29424 25536
rect 0 25168 800 25288
rect 34237 25258 34303 25261
rect 35200 25258 36000 25288
rect 34237 25256 36000 25258
rect 34237 25200 34242 25256
rect 34298 25200 36000 25256
rect 34237 25198 36000 25200
rect 34237 25195 34303 25198
rect 35200 25168 36000 25198
rect 12208 25056 12528 25057
rect 12208 24992 12216 25056
rect 12280 24992 12296 25056
rect 12360 24992 12376 25056
rect 12440 24992 12456 25056
rect 12520 24992 12528 25056
rect 12208 24991 12528 24992
rect 23472 25056 23792 25057
rect 23472 24992 23480 25056
rect 23544 24992 23560 25056
rect 23624 24992 23640 25056
rect 23704 24992 23720 25056
rect 23784 24992 23792 25056
rect 23472 24991 23792 24992
rect 0 24578 800 24608
rect 1485 24578 1551 24581
rect 0 24576 1551 24578
rect 0 24520 1490 24576
rect 1546 24520 1551 24576
rect 0 24518 1551 24520
rect 0 24488 800 24518
rect 1485 24515 1551 24518
rect 34237 24578 34303 24581
rect 35200 24578 36000 24608
rect 34237 24576 36000 24578
rect 34237 24520 34242 24576
rect 34298 24520 36000 24576
rect 34237 24518 36000 24520
rect 34237 24515 34303 24518
rect 6576 24512 6896 24513
rect 6576 24448 6584 24512
rect 6648 24448 6664 24512
rect 6728 24448 6744 24512
rect 6808 24448 6824 24512
rect 6888 24448 6896 24512
rect 6576 24447 6896 24448
rect 17840 24512 18160 24513
rect 17840 24448 17848 24512
rect 17912 24448 17928 24512
rect 17992 24448 18008 24512
rect 18072 24448 18088 24512
rect 18152 24448 18160 24512
rect 17840 24447 18160 24448
rect 29104 24512 29424 24513
rect 29104 24448 29112 24512
rect 29176 24448 29192 24512
rect 29256 24448 29272 24512
rect 29336 24448 29352 24512
rect 29416 24448 29424 24512
rect 35200 24488 36000 24518
rect 29104 24447 29424 24448
rect 12208 23968 12528 23969
rect 0 23898 800 23928
rect 12208 23904 12216 23968
rect 12280 23904 12296 23968
rect 12360 23904 12376 23968
rect 12440 23904 12456 23968
rect 12520 23904 12528 23968
rect 12208 23903 12528 23904
rect 23472 23968 23792 23969
rect 23472 23904 23480 23968
rect 23544 23904 23560 23968
rect 23624 23904 23640 23968
rect 23704 23904 23720 23968
rect 23784 23904 23792 23968
rect 23472 23903 23792 23904
rect 1485 23898 1551 23901
rect 0 23896 1551 23898
rect 0 23840 1490 23896
rect 1546 23840 1551 23896
rect 0 23838 1551 23840
rect 0 23808 800 23838
rect 1485 23835 1551 23838
rect 34237 23898 34303 23901
rect 35200 23898 36000 23928
rect 34237 23896 36000 23898
rect 34237 23840 34242 23896
rect 34298 23840 36000 23896
rect 34237 23838 36000 23840
rect 34237 23835 34303 23838
rect 35200 23808 36000 23838
rect 6576 23424 6896 23425
rect 6576 23360 6584 23424
rect 6648 23360 6664 23424
rect 6728 23360 6744 23424
rect 6808 23360 6824 23424
rect 6888 23360 6896 23424
rect 6576 23359 6896 23360
rect 17840 23424 18160 23425
rect 17840 23360 17848 23424
rect 17912 23360 17928 23424
rect 17992 23360 18008 23424
rect 18072 23360 18088 23424
rect 18152 23360 18160 23424
rect 17840 23359 18160 23360
rect 29104 23424 29424 23425
rect 29104 23360 29112 23424
rect 29176 23360 29192 23424
rect 29256 23360 29272 23424
rect 29336 23360 29352 23424
rect 29416 23360 29424 23424
rect 29104 23359 29424 23360
rect 0 23218 800 23248
rect 1485 23218 1551 23221
rect 0 23216 1551 23218
rect 0 23160 1490 23216
rect 1546 23160 1551 23216
rect 0 23158 1551 23160
rect 0 23128 800 23158
rect 1485 23155 1551 23158
rect 34237 23218 34303 23221
rect 35200 23218 36000 23248
rect 34237 23216 36000 23218
rect 34237 23160 34242 23216
rect 34298 23160 36000 23216
rect 34237 23158 36000 23160
rect 34237 23155 34303 23158
rect 35200 23128 36000 23158
rect 12208 22880 12528 22881
rect 12208 22816 12216 22880
rect 12280 22816 12296 22880
rect 12360 22816 12376 22880
rect 12440 22816 12456 22880
rect 12520 22816 12528 22880
rect 12208 22815 12528 22816
rect 23472 22880 23792 22881
rect 23472 22816 23480 22880
rect 23544 22816 23560 22880
rect 23624 22816 23640 22880
rect 23704 22816 23720 22880
rect 23784 22816 23792 22880
rect 23472 22815 23792 22816
rect 0 22538 800 22568
rect 1485 22538 1551 22541
rect 0 22536 1551 22538
rect 0 22480 1490 22536
rect 1546 22480 1551 22536
rect 0 22478 1551 22480
rect 0 22448 800 22478
rect 1485 22475 1551 22478
rect 34329 22538 34395 22541
rect 35200 22538 36000 22568
rect 34329 22536 36000 22538
rect 34329 22480 34334 22536
rect 34390 22480 36000 22536
rect 34329 22478 36000 22480
rect 34329 22475 34395 22478
rect 35200 22448 36000 22478
rect 6576 22336 6896 22337
rect 6576 22272 6584 22336
rect 6648 22272 6664 22336
rect 6728 22272 6744 22336
rect 6808 22272 6824 22336
rect 6888 22272 6896 22336
rect 6576 22271 6896 22272
rect 17840 22336 18160 22337
rect 17840 22272 17848 22336
rect 17912 22272 17928 22336
rect 17992 22272 18008 22336
rect 18072 22272 18088 22336
rect 18152 22272 18160 22336
rect 17840 22271 18160 22272
rect 29104 22336 29424 22337
rect 29104 22272 29112 22336
rect 29176 22272 29192 22336
rect 29256 22272 29272 22336
rect 29336 22272 29352 22336
rect 29416 22272 29424 22336
rect 29104 22271 29424 22272
rect 12208 21792 12528 21793
rect 12208 21728 12216 21792
rect 12280 21728 12296 21792
rect 12360 21728 12376 21792
rect 12440 21728 12456 21792
rect 12520 21728 12528 21792
rect 12208 21727 12528 21728
rect 23472 21792 23792 21793
rect 23472 21728 23480 21792
rect 23544 21728 23560 21792
rect 23624 21728 23640 21792
rect 23704 21728 23720 21792
rect 23784 21728 23792 21792
rect 23472 21727 23792 21728
rect 6576 21248 6896 21249
rect 0 21178 800 21208
rect 6576 21184 6584 21248
rect 6648 21184 6664 21248
rect 6728 21184 6744 21248
rect 6808 21184 6824 21248
rect 6888 21184 6896 21248
rect 6576 21183 6896 21184
rect 17840 21248 18160 21249
rect 17840 21184 17848 21248
rect 17912 21184 17928 21248
rect 17992 21184 18008 21248
rect 18072 21184 18088 21248
rect 18152 21184 18160 21248
rect 17840 21183 18160 21184
rect 29104 21248 29424 21249
rect 29104 21184 29112 21248
rect 29176 21184 29192 21248
rect 29256 21184 29272 21248
rect 29336 21184 29352 21248
rect 29416 21184 29424 21248
rect 29104 21183 29424 21184
rect 1485 21178 1551 21181
rect 0 21176 1551 21178
rect 0 21120 1490 21176
rect 1546 21120 1551 21176
rect 0 21118 1551 21120
rect 0 21088 800 21118
rect 1485 21115 1551 21118
rect 34329 21178 34395 21181
rect 35200 21178 36000 21208
rect 34329 21176 36000 21178
rect 34329 21120 34334 21176
rect 34390 21120 36000 21176
rect 34329 21118 36000 21120
rect 34329 21115 34395 21118
rect 35200 21088 36000 21118
rect 12208 20704 12528 20705
rect 12208 20640 12216 20704
rect 12280 20640 12296 20704
rect 12360 20640 12376 20704
rect 12440 20640 12456 20704
rect 12520 20640 12528 20704
rect 12208 20639 12528 20640
rect 23472 20704 23792 20705
rect 23472 20640 23480 20704
rect 23544 20640 23560 20704
rect 23624 20640 23640 20704
rect 23704 20640 23720 20704
rect 23784 20640 23792 20704
rect 23472 20639 23792 20640
rect 0 20408 800 20528
rect 33501 20498 33567 20501
rect 35200 20498 36000 20528
rect 33501 20496 36000 20498
rect 33501 20440 33506 20496
rect 33562 20440 36000 20496
rect 33501 20438 36000 20440
rect 33501 20435 33567 20438
rect 35200 20408 36000 20438
rect 6576 20160 6896 20161
rect 6576 20096 6584 20160
rect 6648 20096 6664 20160
rect 6728 20096 6744 20160
rect 6808 20096 6824 20160
rect 6888 20096 6896 20160
rect 6576 20095 6896 20096
rect 17840 20160 18160 20161
rect 17840 20096 17848 20160
rect 17912 20096 17928 20160
rect 17992 20096 18008 20160
rect 18072 20096 18088 20160
rect 18152 20096 18160 20160
rect 17840 20095 18160 20096
rect 29104 20160 29424 20161
rect 29104 20096 29112 20160
rect 29176 20096 29192 20160
rect 29256 20096 29272 20160
rect 29336 20096 29352 20160
rect 29416 20096 29424 20160
rect 29104 20095 29424 20096
rect 0 19818 800 19848
rect 1393 19818 1459 19821
rect 0 19816 1459 19818
rect 0 19760 1398 19816
rect 1454 19760 1459 19816
rect 0 19758 1459 19760
rect 0 19728 800 19758
rect 1393 19755 1459 19758
rect 34329 19818 34395 19821
rect 35200 19818 36000 19848
rect 34329 19816 36000 19818
rect 34329 19760 34334 19816
rect 34390 19760 36000 19816
rect 34329 19758 36000 19760
rect 34329 19755 34395 19758
rect 35200 19728 36000 19758
rect 12208 19616 12528 19617
rect 12208 19552 12216 19616
rect 12280 19552 12296 19616
rect 12360 19552 12376 19616
rect 12440 19552 12456 19616
rect 12520 19552 12528 19616
rect 12208 19551 12528 19552
rect 23472 19616 23792 19617
rect 23472 19552 23480 19616
rect 23544 19552 23560 19616
rect 23624 19552 23640 19616
rect 23704 19552 23720 19616
rect 23784 19552 23792 19616
rect 23472 19551 23792 19552
rect 0 19138 800 19168
rect 1393 19138 1459 19141
rect 0 19136 1459 19138
rect 0 19080 1398 19136
rect 1454 19080 1459 19136
rect 0 19078 1459 19080
rect 0 19048 800 19078
rect 1393 19075 1459 19078
rect 34329 19138 34395 19141
rect 35200 19138 36000 19168
rect 34329 19136 36000 19138
rect 34329 19080 34334 19136
rect 34390 19080 36000 19136
rect 34329 19078 36000 19080
rect 34329 19075 34395 19078
rect 6576 19072 6896 19073
rect 6576 19008 6584 19072
rect 6648 19008 6664 19072
rect 6728 19008 6744 19072
rect 6808 19008 6824 19072
rect 6888 19008 6896 19072
rect 6576 19007 6896 19008
rect 17840 19072 18160 19073
rect 17840 19008 17848 19072
rect 17912 19008 17928 19072
rect 17992 19008 18008 19072
rect 18072 19008 18088 19072
rect 18152 19008 18160 19072
rect 17840 19007 18160 19008
rect 29104 19072 29424 19073
rect 29104 19008 29112 19072
rect 29176 19008 29192 19072
rect 29256 19008 29272 19072
rect 29336 19008 29352 19072
rect 29416 19008 29424 19072
rect 35200 19048 36000 19078
rect 29104 19007 29424 19008
rect 12208 18528 12528 18529
rect 0 18458 800 18488
rect 12208 18464 12216 18528
rect 12280 18464 12296 18528
rect 12360 18464 12376 18528
rect 12440 18464 12456 18528
rect 12520 18464 12528 18528
rect 12208 18463 12528 18464
rect 23472 18528 23792 18529
rect 23472 18464 23480 18528
rect 23544 18464 23560 18528
rect 23624 18464 23640 18528
rect 23704 18464 23720 18528
rect 23784 18464 23792 18528
rect 23472 18463 23792 18464
rect 2129 18458 2195 18461
rect 0 18456 2195 18458
rect 0 18400 2134 18456
rect 2190 18400 2195 18456
rect 0 18398 2195 18400
rect 0 18368 800 18398
rect 2129 18395 2195 18398
rect 34329 18458 34395 18461
rect 35200 18458 36000 18488
rect 34329 18456 36000 18458
rect 34329 18400 34334 18456
rect 34390 18400 36000 18456
rect 34329 18398 36000 18400
rect 34329 18395 34395 18398
rect 35200 18368 36000 18398
rect 6576 17984 6896 17985
rect 6576 17920 6584 17984
rect 6648 17920 6664 17984
rect 6728 17920 6744 17984
rect 6808 17920 6824 17984
rect 6888 17920 6896 17984
rect 6576 17919 6896 17920
rect 17840 17984 18160 17985
rect 17840 17920 17848 17984
rect 17912 17920 17928 17984
rect 17992 17920 18008 17984
rect 18072 17920 18088 17984
rect 18152 17920 18160 17984
rect 17840 17919 18160 17920
rect 29104 17984 29424 17985
rect 29104 17920 29112 17984
rect 29176 17920 29192 17984
rect 29256 17920 29272 17984
rect 29336 17920 29352 17984
rect 29416 17920 29424 17984
rect 29104 17919 29424 17920
rect 0 17778 800 17808
rect 1485 17778 1551 17781
rect 0 17776 1551 17778
rect 0 17720 1490 17776
rect 1546 17720 1551 17776
rect 0 17718 1551 17720
rect 0 17688 800 17718
rect 1485 17715 1551 17718
rect 34237 17778 34303 17781
rect 35200 17778 36000 17808
rect 34237 17776 36000 17778
rect 34237 17720 34242 17776
rect 34298 17720 36000 17776
rect 34237 17718 36000 17720
rect 34237 17715 34303 17718
rect 35200 17688 36000 17718
rect 12208 17440 12528 17441
rect 12208 17376 12216 17440
rect 12280 17376 12296 17440
rect 12360 17376 12376 17440
rect 12440 17376 12456 17440
rect 12520 17376 12528 17440
rect 12208 17375 12528 17376
rect 23472 17440 23792 17441
rect 23472 17376 23480 17440
rect 23544 17376 23560 17440
rect 23624 17376 23640 17440
rect 23704 17376 23720 17440
rect 23784 17376 23792 17440
rect 23472 17375 23792 17376
rect 0 17098 800 17128
rect 1485 17098 1551 17101
rect 0 17096 1551 17098
rect 0 17040 1490 17096
rect 1546 17040 1551 17096
rect 0 17038 1551 17040
rect 0 17008 800 17038
rect 1485 17035 1551 17038
rect 34237 17098 34303 17101
rect 35200 17098 36000 17128
rect 34237 17096 36000 17098
rect 34237 17040 34242 17096
rect 34298 17040 36000 17096
rect 34237 17038 36000 17040
rect 34237 17035 34303 17038
rect 35200 17008 36000 17038
rect 6576 16896 6896 16897
rect 6576 16832 6584 16896
rect 6648 16832 6664 16896
rect 6728 16832 6744 16896
rect 6808 16832 6824 16896
rect 6888 16832 6896 16896
rect 6576 16831 6896 16832
rect 17840 16896 18160 16897
rect 17840 16832 17848 16896
rect 17912 16832 17928 16896
rect 17992 16832 18008 16896
rect 18072 16832 18088 16896
rect 18152 16832 18160 16896
rect 17840 16831 18160 16832
rect 29104 16896 29424 16897
rect 29104 16832 29112 16896
rect 29176 16832 29192 16896
rect 29256 16832 29272 16896
rect 29336 16832 29352 16896
rect 29416 16832 29424 16896
rect 29104 16831 29424 16832
rect 12208 16352 12528 16353
rect 12208 16288 12216 16352
rect 12280 16288 12296 16352
rect 12360 16288 12376 16352
rect 12440 16288 12456 16352
rect 12520 16288 12528 16352
rect 12208 16287 12528 16288
rect 23472 16352 23792 16353
rect 23472 16288 23480 16352
rect 23544 16288 23560 16352
rect 23624 16288 23640 16352
rect 23704 16288 23720 16352
rect 23784 16288 23792 16352
rect 23472 16287 23792 16288
rect 6576 15808 6896 15809
rect 0 15738 800 15768
rect 6576 15744 6584 15808
rect 6648 15744 6664 15808
rect 6728 15744 6744 15808
rect 6808 15744 6824 15808
rect 6888 15744 6896 15808
rect 6576 15743 6896 15744
rect 17840 15808 18160 15809
rect 17840 15744 17848 15808
rect 17912 15744 17928 15808
rect 17992 15744 18008 15808
rect 18072 15744 18088 15808
rect 18152 15744 18160 15808
rect 17840 15743 18160 15744
rect 29104 15808 29424 15809
rect 29104 15744 29112 15808
rect 29176 15744 29192 15808
rect 29256 15744 29272 15808
rect 29336 15744 29352 15808
rect 29416 15744 29424 15808
rect 29104 15743 29424 15744
rect 1485 15738 1551 15741
rect 0 15736 1551 15738
rect 0 15680 1490 15736
rect 1546 15680 1551 15736
rect 0 15678 1551 15680
rect 0 15648 800 15678
rect 1485 15675 1551 15678
rect 34329 15738 34395 15741
rect 35200 15738 36000 15768
rect 34329 15736 36000 15738
rect 34329 15680 34334 15736
rect 34390 15680 36000 15736
rect 34329 15678 36000 15680
rect 34329 15675 34395 15678
rect 35200 15648 36000 15678
rect 12208 15264 12528 15265
rect 12208 15200 12216 15264
rect 12280 15200 12296 15264
rect 12360 15200 12376 15264
rect 12440 15200 12456 15264
rect 12520 15200 12528 15264
rect 12208 15199 12528 15200
rect 23472 15264 23792 15265
rect 23472 15200 23480 15264
rect 23544 15200 23560 15264
rect 23624 15200 23640 15264
rect 23704 15200 23720 15264
rect 23784 15200 23792 15264
rect 23472 15199 23792 15200
rect 0 15058 800 15088
rect 1393 15058 1459 15061
rect 0 15056 1459 15058
rect 0 15000 1398 15056
rect 1454 15000 1459 15056
rect 0 14998 1459 15000
rect 0 14968 800 14998
rect 1393 14995 1459 14998
rect 34237 15058 34303 15061
rect 35200 15058 36000 15088
rect 34237 15056 36000 15058
rect 34237 15000 34242 15056
rect 34298 15000 36000 15056
rect 34237 14998 36000 15000
rect 34237 14995 34303 14998
rect 35200 14968 36000 14998
rect 6576 14720 6896 14721
rect 6576 14656 6584 14720
rect 6648 14656 6664 14720
rect 6728 14656 6744 14720
rect 6808 14656 6824 14720
rect 6888 14656 6896 14720
rect 6576 14655 6896 14656
rect 17840 14720 18160 14721
rect 17840 14656 17848 14720
rect 17912 14656 17928 14720
rect 17992 14656 18008 14720
rect 18072 14656 18088 14720
rect 18152 14656 18160 14720
rect 17840 14655 18160 14656
rect 29104 14720 29424 14721
rect 29104 14656 29112 14720
rect 29176 14656 29192 14720
rect 29256 14656 29272 14720
rect 29336 14656 29352 14720
rect 29416 14656 29424 14720
rect 29104 14655 29424 14656
rect 0 14378 800 14408
rect 1485 14378 1551 14381
rect 0 14376 1551 14378
rect 0 14320 1490 14376
rect 1546 14320 1551 14376
rect 0 14318 1551 14320
rect 0 14288 800 14318
rect 1485 14315 1551 14318
rect 34329 14378 34395 14381
rect 35200 14378 36000 14408
rect 34329 14376 36000 14378
rect 34329 14320 34334 14376
rect 34390 14320 36000 14376
rect 34329 14318 36000 14320
rect 34329 14315 34395 14318
rect 35200 14288 36000 14318
rect 12208 14176 12528 14177
rect 12208 14112 12216 14176
rect 12280 14112 12296 14176
rect 12360 14112 12376 14176
rect 12440 14112 12456 14176
rect 12520 14112 12528 14176
rect 12208 14111 12528 14112
rect 23472 14176 23792 14177
rect 23472 14112 23480 14176
rect 23544 14112 23560 14176
rect 23624 14112 23640 14176
rect 23704 14112 23720 14176
rect 23784 14112 23792 14176
rect 23472 14111 23792 14112
rect 0 13608 800 13728
rect 34329 13698 34395 13701
rect 35200 13698 36000 13728
rect 34329 13696 36000 13698
rect 34329 13640 34334 13696
rect 34390 13640 36000 13696
rect 34329 13638 36000 13640
rect 34329 13635 34395 13638
rect 6576 13632 6896 13633
rect 6576 13568 6584 13632
rect 6648 13568 6664 13632
rect 6728 13568 6744 13632
rect 6808 13568 6824 13632
rect 6888 13568 6896 13632
rect 6576 13567 6896 13568
rect 17840 13632 18160 13633
rect 17840 13568 17848 13632
rect 17912 13568 17928 13632
rect 17992 13568 18008 13632
rect 18072 13568 18088 13632
rect 18152 13568 18160 13632
rect 17840 13567 18160 13568
rect 29104 13632 29424 13633
rect 29104 13568 29112 13632
rect 29176 13568 29192 13632
rect 29256 13568 29272 13632
rect 29336 13568 29352 13632
rect 29416 13568 29424 13632
rect 35200 13608 36000 13638
rect 29104 13567 29424 13568
rect 12208 13088 12528 13089
rect 0 13018 800 13048
rect 12208 13024 12216 13088
rect 12280 13024 12296 13088
rect 12360 13024 12376 13088
rect 12440 13024 12456 13088
rect 12520 13024 12528 13088
rect 12208 13023 12528 13024
rect 23472 13088 23792 13089
rect 23472 13024 23480 13088
rect 23544 13024 23560 13088
rect 23624 13024 23640 13088
rect 23704 13024 23720 13088
rect 23784 13024 23792 13088
rect 23472 13023 23792 13024
rect 1669 13018 1735 13021
rect 0 13016 1735 13018
rect 0 12960 1674 13016
rect 1730 12960 1735 13016
rect 0 12958 1735 12960
rect 0 12928 800 12958
rect 1669 12955 1735 12958
rect 34237 13018 34303 13021
rect 35200 13018 36000 13048
rect 34237 13016 36000 13018
rect 34237 12960 34242 13016
rect 34298 12960 36000 13016
rect 34237 12958 36000 12960
rect 34237 12955 34303 12958
rect 35200 12928 36000 12958
rect 6576 12544 6896 12545
rect 6576 12480 6584 12544
rect 6648 12480 6664 12544
rect 6728 12480 6744 12544
rect 6808 12480 6824 12544
rect 6888 12480 6896 12544
rect 6576 12479 6896 12480
rect 17840 12544 18160 12545
rect 17840 12480 17848 12544
rect 17912 12480 17928 12544
rect 17992 12480 18008 12544
rect 18072 12480 18088 12544
rect 18152 12480 18160 12544
rect 17840 12479 18160 12480
rect 29104 12544 29424 12545
rect 29104 12480 29112 12544
rect 29176 12480 29192 12544
rect 29256 12480 29272 12544
rect 29336 12480 29352 12544
rect 29416 12480 29424 12544
rect 29104 12479 29424 12480
rect 0 12338 800 12368
rect 1485 12338 1551 12341
rect 0 12336 1551 12338
rect 0 12280 1490 12336
rect 1546 12280 1551 12336
rect 0 12278 1551 12280
rect 0 12248 800 12278
rect 1485 12275 1551 12278
rect 34237 12338 34303 12341
rect 35200 12338 36000 12368
rect 34237 12336 36000 12338
rect 34237 12280 34242 12336
rect 34298 12280 36000 12336
rect 34237 12278 36000 12280
rect 34237 12275 34303 12278
rect 35200 12248 36000 12278
rect 12208 12000 12528 12001
rect 12208 11936 12216 12000
rect 12280 11936 12296 12000
rect 12360 11936 12376 12000
rect 12440 11936 12456 12000
rect 12520 11936 12528 12000
rect 12208 11935 12528 11936
rect 23472 12000 23792 12001
rect 23472 11936 23480 12000
rect 23544 11936 23560 12000
rect 23624 11936 23640 12000
rect 23704 11936 23720 12000
rect 23784 11936 23792 12000
rect 23472 11935 23792 11936
rect 0 11658 800 11688
rect 1393 11658 1459 11661
rect 0 11656 1459 11658
rect 0 11600 1398 11656
rect 1454 11600 1459 11656
rect 0 11598 1459 11600
rect 0 11568 800 11598
rect 1393 11595 1459 11598
rect 34237 11658 34303 11661
rect 35200 11658 36000 11688
rect 34237 11656 36000 11658
rect 34237 11600 34242 11656
rect 34298 11600 36000 11656
rect 34237 11598 36000 11600
rect 34237 11595 34303 11598
rect 35200 11568 36000 11598
rect 6576 11456 6896 11457
rect 6576 11392 6584 11456
rect 6648 11392 6664 11456
rect 6728 11392 6744 11456
rect 6808 11392 6824 11456
rect 6888 11392 6896 11456
rect 6576 11391 6896 11392
rect 17840 11456 18160 11457
rect 17840 11392 17848 11456
rect 17912 11392 17928 11456
rect 17992 11392 18008 11456
rect 18072 11392 18088 11456
rect 18152 11392 18160 11456
rect 17840 11391 18160 11392
rect 29104 11456 29424 11457
rect 29104 11392 29112 11456
rect 29176 11392 29192 11456
rect 29256 11392 29272 11456
rect 29336 11392 29352 11456
rect 29416 11392 29424 11456
rect 29104 11391 29424 11392
rect 12208 10912 12528 10913
rect 12208 10848 12216 10912
rect 12280 10848 12296 10912
rect 12360 10848 12376 10912
rect 12440 10848 12456 10912
rect 12520 10848 12528 10912
rect 12208 10847 12528 10848
rect 23472 10912 23792 10913
rect 23472 10848 23480 10912
rect 23544 10848 23560 10912
rect 23624 10848 23640 10912
rect 23704 10848 23720 10912
rect 23784 10848 23792 10912
rect 23472 10847 23792 10848
rect 6576 10368 6896 10369
rect 0 10298 800 10328
rect 6576 10304 6584 10368
rect 6648 10304 6664 10368
rect 6728 10304 6744 10368
rect 6808 10304 6824 10368
rect 6888 10304 6896 10368
rect 6576 10303 6896 10304
rect 17840 10368 18160 10369
rect 17840 10304 17848 10368
rect 17912 10304 17928 10368
rect 17992 10304 18008 10368
rect 18072 10304 18088 10368
rect 18152 10304 18160 10368
rect 17840 10303 18160 10304
rect 29104 10368 29424 10369
rect 29104 10304 29112 10368
rect 29176 10304 29192 10368
rect 29256 10304 29272 10368
rect 29336 10304 29352 10368
rect 29416 10304 29424 10368
rect 29104 10303 29424 10304
rect 1393 10298 1459 10301
rect 0 10296 1459 10298
rect 0 10240 1398 10296
rect 1454 10240 1459 10296
rect 0 10238 1459 10240
rect 0 10208 800 10238
rect 1393 10235 1459 10238
rect 35200 10208 36000 10328
rect 12208 9824 12528 9825
rect 12208 9760 12216 9824
rect 12280 9760 12296 9824
rect 12360 9760 12376 9824
rect 12440 9760 12456 9824
rect 12520 9760 12528 9824
rect 12208 9759 12528 9760
rect 23472 9824 23792 9825
rect 23472 9760 23480 9824
rect 23544 9760 23560 9824
rect 23624 9760 23640 9824
rect 23704 9760 23720 9824
rect 23784 9760 23792 9824
rect 23472 9759 23792 9760
rect 0 9528 800 9648
rect 34329 9618 34395 9621
rect 35200 9618 36000 9648
rect 34329 9616 36000 9618
rect 34329 9560 34334 9616
rect 34390 9560 36000 9616
rect 34329 9558 36000 9560
rect 34329 9555 34395 9558
rect 35200 9528 36000 9558
rect 6576 9280 6896 9281
rect 6576 9216 6584 9280
rect 6648 9216 6664 9280
rect 6728 9216 6744 9280
rect 6808 9216 6824 9280
rect 6888 9216 6896 9280
rect 6576 9215 6896 9216
rect 17840 9280 18160 9281
rect 17840 9216 17848 9280
rect 17912 9216 17928 9280
rect 17992 9216 18008 9280
rect 18072 9216 18088 9280
rect 18152 9216 18160 9280
rect 17840 9215 18160 9216
rect 29104 9280 29424 9281
rect 29104 9216 29112 9280
rect 29176 9216 29192 9280
rect 29256 9216 29272 9280
rect 29336 9216 29352 9280
rect 29416 9216 29424 9280
rect 29104 9215 29424 9216
rect 0 8938 800 8968
rect 1485 8938 1551 8941
rect 0 8936 1551 8938
rect 0 8880 1490 8936
rect 1546 8880 1551 8936
rect 0 8878 1551 8880
rect 0 8848 800 8878
rect 1485 8875 1551 8878
rect 34237 8938 34303 8941
rect 35200 8938 36000 8968
rect 34237 8936 36000 8938
rect 34237 8880 34242 8936
rect 34298 8880 36000 8936
rect 34237 8878 36000 8880
rect 34237 8875 34303 8878
rect 35200 8848 36000 8878
rect 12208 8736 12528 8737
rect 12208 8672 12216 8736
rect 12280 8672 12296 8736
rect 12360 8672 12376 8736
rect 12440 8672 12456 8736
rect 12520 8672 12528 8736
rect 12208 8671 12528 8672
rect 23472 8736 23792 8737
rect 23472 8672 23480 8736
rect 23544 8672 23560 8736
rect 23624 8672 23640 8736
rect 23704 8672 23720 8736
rect 23784 8672 23792 8736
rect 23472 8671 23792 8672
rect 0 8168 800 8288
rect 34237 8258 34303 8261
rect 35200 8258 36000 8288
rect 34237 8256 36000 8258
rect 34237 8200 34242 8256
rect 34298 8200 36000 8256
rect 34237 8198 36000 8200
rect 34237 8195 34303 8198
rect 6576 8192 6896 8193
rect 6576 8128 6584 8192
rect 6648 8128 6664 8192
rect 6728 8128 6744 8192
rect 6808 8128 6824 8192
rect 6888 8128 6896 8192
rect 6576 8127 6896 8128
rect 17840 8192 18160 8193
rect 17840 8128 17848 8192
rect 17912 8128 17928 8192
rect 17992 8128 18008 8192
rect 18072 8128 18088 8192
rect 18152 8128 18160 8192
rect 17840 8127 18160 8128
rect 29104 8192 29424 8193
rect 29104 8128 29112 8192
rect 29176 8128 29192 8192
rect 29256 8128 29272 8192
rect 29336 8128 29352 8192
rect 29416 8128 29424 8192
rect 35200 8168 36000 8198
rect 29104 8127 29424 8128
rect 12208 7648 12528 7649
rect 0 7578 800 7608
rect 12208 7584 12216 7648
rect 12280 7584 12296 7648
rect 12360 7584 12376 7648
rect 12440 7584 12456 7648
rect 12520 7584 12528 7648
rect 12208 7583 12528 7584
rect 23472 7648 23792 7649
rect 23472 7584 23480 7648
rect 23544 7584 23560 7648
rect 23624 7584 23640 7648
rect 23704 7584 23720 7648
rect 23784 7584 23792 7648
rect 23472 7583 23792 7584
rect 1485 7578 1551 7581
rect 0 7576 1551 7578
rect 0 7520 1490 7576
rect 1546 7520 1551 7576
rect 0 7518 1551 7520
rect 0 7488 800 7518
rect 1485 7515 1551 7518
rect 34237 7578 34303 7581
rect 35200 7578 36000 7608
rect 34237 7576 36000 7578
rect 34237 7520 34242 7576
rect 34298 7520 36000 7576
rect 34237 7518 36000 7520
rect 34237 7515 34303 7518
rect 35200 7488 36000 7518
rect 6576 7104 6896 7105
rect 6576 7040 6584 7104
rect 6648 7040 6664 7104
rect 6728 7040 6744 7104
rect 6808 7040 6824 7104
rect 6888 7040 6896 7104
rect 6576 7039 6896 7040
rect 17840 7104 18160 7105
rect 17840 7040 17848 7104
rect 17912 7040 17928 7104
rect 17992 7040 18008 7104
rect 18072 7040 18088 7104
rect 18152 7040 18160 7104
rect 17840 7039 18160 7040
rect 29104 7104 29424 7105
rect 29104 7040 29112 7104
rect 29176 7040 29192 7104
rect 29256 7040 29272 7104
rect 29336 7040 29352 7104
rect 29416 7040 29424 7104
rect 29104 7039 29424 7040
rect 0 6898 800 6928
rect 1485 6898 1551 6901
rect 0 6896 1551 6898
rect 0 6840 1490 6896
rect 1546 6840 1551 6896
rect 0 6838 1551 6840
rect 0 6808 800 6838
rect 1485 6835 1551 6838
rect 34237 6898 34303 6901
rect 35200 6898 36000 6928
rect 34237 6896 36000 6898
rect 34237 6840 34242 6896
rect 34298 6840 36000 6896
rect 34237 6838 36000 6840
rect 34237 6835 34303 6838
rect 35200 6808 36000 6838
rect 12208 6560 12528 6561
rect 12208 6496 12216 6560
rect 12280 6496 12296 6560
rect 12360 6496 12376 6560
rect 12440 6496 12456 6560
rect 12520 6496 12528 6560
rect 12208 6495 12528 6496
rect 23472 6560 23792 6561
rect 23472 6496 23480 6560
rect 23544 6496 23560 6560
rect 23624 6496 23640 6560
rect 23704 6496 23720 6560
rect 23784 6496 23792 6560
rect 23472 6495 23792 6496
rect 0 6218 800 6248
rect 1485 6218 1551 6221
rect 0 6216 1551 6218
rect 0 6160 1490 6216
rect 1546 6160 1551 6216
rect 0 6158 1551 6160
rect 0 6128 800 6158
rect 1485 6155 1551 6158
rect 34237 6218 34303 6221
rect 35200 6218 36000 6248
rect 34237 6216 36000 6218
rect 34237 6160 34242 6216
rect 34298 6160 36000 6216
rect 34237 6158 36000 6160
rect 34237 6155 34303 6158
rect 35200 6128 36000 6158
rect 6576 6016 6896 6017
rect 6576 5952 6584 6016
rect 6648 5952 6664 6016
rect 6728 5952 6744 6016
rect 6808 5952 6824 6016
rect 6888 5952 6896 6016
rect 6576 5951 6896 5952
rect 17840 6016 18160 6017
rect 17840 5952 17848 6016
rect 17912 5952 17928 6016
rect 17992 5952 18008 6016
rect 18072 5952 18088 6016
rect 18152 5952 18160 6016
rect 17840 5951 18160 5952
rect 29104 6016 29424 6017
rect 29104 5952 29112 6016
rect 29176 5952 29192 6016
rect 29256 5952 29272 6016
rect 29336 5952 29352 6016
rect 29416 5952 29424 6016
rect 29104 5951 29424 5952
rect 12208 5472 12528 5473
rect 12208 5408 12216 5472
rect 12280 5408 12296 5472
rect 12360 5408 12376 5472
rect 12440 5408 12456 5472
rect 12520 5408 12528 5472
rect 12208 5407 12528 5408
rect 23472 5472 23792 5473
rect 23472 5408 23480 5472
rect 23544 5408 23560 5472
rect 23624 5408 23640 5472
rect 23704 5408 23720 5472
rect 23784 5408 23792 5472
rect 23472 5407 23792 5408
rect 6576 4928 6896 4929
rect 0 4858 800 4888
rect 6576 4864 6584 4928
rect 6648 4864 6664 4928
rect 6728 4864 6744 4928
rect 6808 4864 6824 4928
rect 6888 4864 6896 4928
rect 6576 4863 6896 4864
rect 17840 4928 18160 4929
rect 17840 4864 17848 4928
rect 17912 4864 17928 4928
rect 17992 4864 18008 4928
rect 18072 4864 18088 4928
rect 18152 4864 18160 4928
rect 17840 4863 18160 4864
rect 29104 4928 29424 4929
rect 29104 4864 29112 4928
rect 29176 4864 29192 4928
rect 29256 4864 29272 4928
rect 29336 4864 29352 4928
rect 29416 4864 29424 4928
rect 29104 4863 29424 4864
rect 1485 4858 1551 4861
rect 0 4856 1551 4858
rect 0 4800 1490 4856
rect 1546 4800 1551 4856
rect 0 4798 1551 4800
rect 0 4768 800 4798
rect 1485 4795 1551 4798
rect 34329 4858 34395 4861
rect 35200 4858 36000 4888
rect 34329 4856 36000 4858
rect 34329 4800 34334 4856
rect 34390 4800 36000 4856
rect 34329 4798 36000 4800
rect 34329 4795 34395 4798
rect 35200 4768 36000 4798
rect 12208 4384 12528 4385
rect 12208 4320 12216 4384
rect 12280 4320 12296 4384
rect 12360 4320 12376 4384
rect 12440 4320 12456 4384
rect 12520 4320 12528 4384
rect 12208 4319 12528 4320
rect 23472 4384 23792 4385
rect 23472 4320 23480 4384
rect 23544 4320 23560 4384
rect 23624 4320 23640 4384
rect 23704 4320 23720 4384
rect 23784 4320 23792 4384
rect 23472 4319 23792 4320
rect 0 4088 800 4208
rect 34237 4178 34303 4181
rect 35200 4178 36000 4208
rect 34237 4176 36000 4178
rect 34237 4120 34242 4176
rect 34298 4120 36000 4176
rect 34237 4118 36000 4120
rect 34237 4115 34303 4118
rect 35200 4088 36000 4118
rect 6576 3840 6896 3841
rect 6576 3776 6584 3840
rect 6648 3776 6664 3840
rect 6728 3776 6744 3840
rect 6808 3776 6824 3840
rect 6888 3776 6896 3840
rect 6576 3775 6896 3776
rect 17840 3840 18160 3841
rect 17840 3776 17848 3840
rect 17912 3776 17928 3840
rect 17992 3776 18008 3840
rect 18072 3776 18088 3840
rect 18152 3776 18160 3840
rect 17840 3775 18160 3776
rect 29104 3840 29424 3841
rect 29104 3776 29112 3840
rect 29176 3776 29192 3840
rect 29256 3776 29272 3840
rect 29336 3776 29352 3840
rect 29416 3776 29424 3840
rect 29104 3775 29424 3776
rect 0 3408 800 3528
rect 19057 3498 19123 3501
rect 32397 3498 32463 3501
rect 19057 3496 32463 3498
rect 19057 3440 19062 3496
rect 19118 3440 32402 3496
rect 32458 3440 32463 3496
rect 19057 3438 32463 3440
rect 19057 3435 19123 3438
rect 32397 3435 32463 3438
rect 35200 3408 36000 3528
rect 12208 3296 12528 3297
rect 12208 3232 12216 3296
rect 12280 3232 12296 3296
rect 12360 3232 12376 3296
rect 12440 3232 12456 3296
rect 12520 3232 12528 3296
rect 12208 3231 12528 3232
rect 23472 3296 23792 3297
rect 23472 3232 23480 3296
rect 23544 3232 23560 3296
rect 23624 3232 23640 3296
rect 23704 3232 23720 3296
rect 23784 3232 23792 3296
rect 23472 3231 23792 3232
rect 0 2818 800 2848
rect 1393 2818 1459 2821
rect 0 2816 1459 2818
rect 0 2760 1398 2816
rect 1454 2760 1459 2816
rect 0 2758 1459 2760
rect 0 2728 800 2758
rect 1393 2755 1459 2758
rect 34237 2818 34303 2821
rect 35200 2818 36000 2848
rect 34237 2816 36000 2818
rect 34237 2760 34242 2816
rect 34298 2760 36000 2816
rect 34237 2758 36000 2760
rect 34237 2755 34303 2758
rect 6576 2752 6896 2753
rect 6576 2688 6584 2752
rect 6648 2688 6664 2752
rect 6728 2688 6744 2752
rect 6808 2688 6824 2752
rect 6888 2688 6896 2752
rect 6576 2687 6896 2688
rect 17840 2752 18160 2753
rect 17840 2688 17848 2752
rect 17912 2688 17928 2752
rect 17992 2688 18008 2752
rect 18072 2688 18088 2752
rect 18152 2688 18160 2752
rect 17840 2687 18160 2688
rect 29104 2752 29424 2753
rect 29104 2688 29112 2752
rect 29176 2688 29192 2752
rect 29256 2688 29272 2752
rect 29336 2688 29352 2752
rect 29416 2688 29424 2752
rect 35200 2728 36000 2758
rect 29104 2687 29424 2688
rect 12208 2208 12528 2209
rect 0 2138 800 2168
rect 12208 2144 12216 2208
rect 12280 2144 12296 2208
rect 12360 2144 12376 2208
rect 12440 2144 12456 2208
rect 12520 2144 12528 2208
rect 12208 2143 12528 2144
rect 23472 2208 23792 2209
rect 23472 2144 23480 2208
rect 23544 2144 23560 2208
rect 23624 2144 23640 2208
rect 23704 2144 23720 2208
rect 23784 2144 23792 2208
rect 23472 2143 23792 2144
rect 2865 2138 2931 2141
rect 0 2136 2931 2138
rect 0 2080 2870 2136
rect 2926 2080 2931 2136
rect 0 2078 2931 2080
rect 0 2048 800 2078
rect 2865 2075 2931 2078
rect 32581 2138 32647 2141
rect 35200 2138 36000 2168
rect 32581 2136 36000 2138
rect 32581 2080 32586 2136
rect 32642 2080 36000 2136
rect 32581 2078 36000 2080
rect 32581 2075 32647 2078
rect 35200 2048 36000 2078
rect 0 1458 800 1488
rect 2957 1458 3023 1461
rect 0 1456 3023 1458
rect 0 1400 2962 1456
rect 3018 1400 3023 1456
rect 0 1398 3023 1400
rect 0 1368 800 1398
rect 2957 1395 3023 1398
rect 33133 1458 33199 1461
rect 35200 1458 36000 1488
rect 33133 1456 36000 1458
rect 33133 1400 33138 1456
rect 33194 1400 36000 1456
rect 33133 1398 36000 1400
rect 33133 1395 33199 1398
rect 35200 1368 36000 1398
rect 0 778 800 808
rect 2957 778 3023 781
rect 0 776 3023 778
rect 0 720 2962 776
rect 3018 720 3023 776
rect 0 718 3023 720
rect 0 688 800 718
rect 2957 715 3023 718
rect 33869 778 33935 781
rect 35200 778 36000 808
rect 33869 776 36000 778
rect 33869 720 33874 776
rect 33930 720 36000 776
rect 33869 718 36000 720
rect 33869 715 33935 718
rect 35200 688 36000 718
<< via3 >>
rect 12216 33756 12280 33760
rect 12216 33700 12220 33756
rect 12220 33700 12276 33756
rect 12276 33700 12280 33756
rect 12216 33696 12280 33700
rect 12296 33756 12360 33760
rect 12296 33700 12300 33756
rect 12300 33700 12356 33756
rect 12356 33700 12360 33756
rect 12296 33696 12360 33700
rect 12376 33756 12440 33760
rect 12376 33700 12380 33756
rect 12380 33700 12436 33756
rect 12436 33700 12440 33756
rect 12376 33696 12440 33700
rect 12456 33756 12520 33760
rect 12456 33700 12460 33756
rect 12460 33700 12516 33756
rect 12516 33700 12520 33756
rect 12456 33696 12520 33700
rect 23480 33756 23544 33760
rect 23480 33700 23484 33756
rect 23484 33700 23540 33756
rect 23540 33700 23544 33756
rect 23480 33696 23544 33700
rect 23560 33756 23624 33760
rect 23560 33700 23564 33756
rect 23564 33700 23620 33756
rect 23620 33700 23624 33756
rect 23560 33696 23624 33700
rect 23640 33756 23704 33760
rect 23640 33700 23644 33756
rect 23644 33700 23700 33756
rect 23700 33700 23704 33756
rect 23640 33696 23704 33700
rect 23720 33756 23784 33760
rect 23720 33700 23724 33756
rect 23724 33700 23780 33756
rect 23780 33700 23784 33756
rect 23720 33696 23784 33700
rect 6584 33212 6648 33216
rect 6584 33156 6588 33212
rect 6588 33156 6644 33212
rect 6644 33156 6648 33212
rect 6584 33152 6648 33156
rect 6664 33212 6728 33216
rect 6664 33156 6668 33212
rect 6668 33156 6724 33212
rect 6724 33156 6728 33212
rect 6664 33152 6728 33156
rect 6744 33212 6808 33216
rect 6744 33156 6748 33212
rect 6748 33156 6804 33212
rect 6804 33156 6808 33212
rect 6744 33152 6808 33156
rect 6824 33212 6888 33216
rect 6824 33156 6828 33212
rect 6828 33156 6884 33212
rect 6884 33156 6888 33212
rect 6824 33152 6888 33156
rect 17848 33212 17912 33216
rect 17848 33156 17852 33212
rect 17852 33156 17908 33212
rect 17908 33156 17912 33212
rect 17848 33152 17912 33156
rect 17928 33212 17992 33216
rect 17928 33156 17932 33212
rect 17932 33156 17988 33212
rect 17988 33156 17992 33212
rect 17928 33152 17992 33156
rect 18008 33212 18072 33216
rect 18008 33156 18012 33212
rect 18012 33156 18068 33212
rect 18068 33156 18072 33212
rect 18008 33152 18072 33156
rect 18088 33212 18152 33216
rect 18088 33156 18092 33212
rect 18092 33156 18148 33212
rect 18148 33156 18152 33212
rect 18088 33152 18152 33156
rect 29112 33212 29176 33216
rect 29112 33156 29116 33212
rect 29116 33156 29172 33212
rect 29172 33156 29176 33212
rect 29112 33152 29176 33156
rect 29192 33212 29256 33216
rect 29192 33156 29196 33212
rect 29196 33156 29252 33212
rect 29252 33156 29256 33212
rect 29192 33152 29256 33156
rect 29272 33212 29336 33216
rect 29272 33156 29276 33212
rect 29276 33156 29332 33212
rect 29332 33156 29336 33212
rect 29272 33152 29336 33156
rect 29352 33212 29416 33216
rect 29352 33156 29356 33212
rect 29356 33156 29412 33212
rect 29412 33156 29416 33212
rect 29352 33152 29416 33156
rect 12216 32668 12280 32672
rect 12216 32612 12220 32668
rect 12220 32612 12276 32668
rect 12276 32612 12280 32668
rect 12216 32608 12280 32612
rect 12296 32668 12360 32672
rect 12296 32612 12300 32668
rect 12300 32612 12356 32668
rect 12356 32612 12360 32668
rect 12296 32608 12360 32612
rect 12376 32668 12440 32672
rect 12376 32612 12380 32668
rect 12380 32612 12436 32668
rect 12436 32612 12440 32668
rect 12376 32608 12440 32612
rect 12456 32668 12520 32672
rect 12456 32612 12460 32668
rect 12460 32612 12516 32668
rect 12516 32612 12520 32668
rect 12456 32608 12520 32612
rect 23480 32668 23544 32672
rect 23480 32612 23484 32668
rect 23484 32612 23540 32668
rect 23540 32612 23544 32668
rect 23480 32608 23544 32612
rect 23560 32668 23624 32672
rect 23560 32612 23564 32668
rect 23564 32612 23620 32668
rect 23620 32612 23624 32668
rect 23560 32608 23624 32612
rect 23640 32668 23704 32672
rect 23640 32612 23644 32668
rect 23644 32612 23700 32668
rect 23700 32612 23704 32668
rect 23640 32608 23704 32612
rect 23720 32668 23784 32672
rect 23720 32612 23724 32668
rect 23724 32612 23780 32668
rect 23780 32612 23784 32668
rect 23720 32608 23784 32612
rect 6584 32124 6648 32128
rect 6584 32068 6588 32124
rect 6588 32068 6644 32124
rect 6644 32068 6648 32124
rect 6584 32064 6648 32068
rect 6664 32124 6728 32128
rect 6664 32068 6668 32124
rect 6668 32068 6724 32124
rect 6724 32068 6728 32124
rect 6664 32064 6728 32068
rect 6744 32124 6808 32128
rect 6744 32068 6748 32124
rect 6748 32068 6804 32124
rect 6804 32068 6808 32124
rect 6744 32064 6808 32068
rect 6824 32124 6888 32128
rect 6824 32068 6828 32124
rect 6828 32068 6884 32124
rect 6884 32068 6888 32124
rect 6824 32064 6888 32068
rect 17848 32124 17912 32128
rect 17848 32068 17852 32124
rect 17852 32068 17908 32124
rect 17908 32068 17912 32124
rect 17848 32064 17912 32068
rect 17928 32124 17992 32128
rect 17928 32068 17932 32124
rect 17932 32068 17988 32124
rect 17988 32068 17992 32124
rect 17928 32064 17992 32068
rect 18008 32124 18072 32128
rect 18008 32068 18012 32124
rect 18012 32068 18068 32124
rect 18068 32068 18072 32124
rect 18008 32064 18072 32068
rect 18088 32124 18152 32128
rect 18088 32068 18092 32124
rect 18092 32068 18148 32124
rect 18148 32068 18152 32124
rect 18088 32064 18152 32068
rect 29112 32124 29176 32128
rect 29112 32068 29116 32124
rect 29116 32068 29172 32124
rect 29172 32068 29176 32124
rect 29112 32064 29176 32068
rect 29192 32124 29256 32128
rect 29192 32068 29196 32124
rect 29196 32068 29252 32124
rect 29252 32068 29256 32124
rect 29192 32064 29256 32068
rect 29272 32124 29336 32128
rect 29272 32068 29276 32124
rect 29276 32068 29332 32124
rect 29332 32068 29336 32124
rect 29272 32064 29336 32068
rect 29352 32124 29416 32128
rect 29352 32068 29356 32124
rect 29356 32068 29412 32124
rect 29412 32068 29416 32124
rect 29352 32064 29416 32068
rect 12216 31580 12280 31584
rect 12216 31524 12220 31580
rect 12220 31524 12276 31580
rect 12276 31524 12280 31580
rect 12216 31520 12280 31524
rect 12296 31580 12360 31584
rect 12296 31524 12300 31580
rect 12300 31524 12356 31580
rect 12356 31524 12360 31580
rect 12296 31520 12360 31524
rect 12376 31580 12440 31584
rect 12376 31524 12380 31580
rect 12380 31524 12436 31580
rect 12436 31524 12440 31580
rect 12376 31520 12440 31524
rect 12456 31580 12520 31584
rect 12456 31524 12460 31580
rect 12460 31524 12516 31580
rect 12516 31524 12520 31580
rect 12456 31520 12520 31524
rect 23480 31580 23544 31584
rect 23480 31524 23484 31580
rect 23484 31524 23540 31580
rect 23540 31524 23544 31580
rect 23480 31520 23544 31524
rect 23560 31580 23624 31584
rect 23560 31524 23564 31580
rect 23564 31524 23620 31580
rect 23620 31524 23624 31580
rect 23560 31520 23624 31524
rect 23640 31580 23704 31584
rect 23640 31524 23644 31580
rect 23644 31524 23700 31580
rect 23700 31524 23704 31580
rect 23640 31520 23704 31524
rect 23720 31580 23784 31584
rect 23720 31524 23724 31580
rect 23724 31524 23780 31580
rect 23780 31524 23784 31580
rect 23720 31520 23784 31524
rect 6584 31036 6648 31040
rect 6584 30980 6588 31036
rect 6588 30980 6644 31036
rect 6644 30980 6648 31036
rect 6584 30976 6648 30980
rect 6664 31036 6728 31040
rect 6664 30980 6668 31036
rect 6668 30980 6724 31036
rect 6724 30980 6728 31036
rect 6664 30976 6728 30980
rect 6744 31036 6808 31040
rect 6744 30980 6748 31036
rect 6748 30980 6804 31036
rect 6804 30980 6808 31036
rect 6744 30976 6808 30980
rect 6824 31036 6888 31040
rect 6824 30980 6828 31036
rect 6828 30980 6884 31036
rect 6884 30980 6888 31036
rect 6824 30976 6888 30980
rect 17848 31036 17912 31040
rect 17848 30980 17852 31036
rect 17852 30980 17908 31036
rect 17908 30980 17912 31036
rect 17848 30976 17912 30980
rect 17928 31036 17992 31040
rect 17928 30980 17932 31036
rect 17932 30980 17988 31036
rect 17988 30980 17992 31036
rect 17928 30976 17992 30980
rect 18008 31036 18072 31040
rect 18008 30980 18012 31036
rect 18012 30980 18068 31036
rect 18068 30980 18072 31036
rect 18008 30976 18072 30980
rect 18088 31036 18152 31040
rect 18088 30980 18092 31036
rect 18092 30980 18148 31036
rect 18148 30980 18152 31036
rect 18088 30976 18152 30980
rect 29112 31036 29176 31040
rect 29112 30980 29116 31036
rect 29116 30980 29172 31036
rect 29172 30980 29176 31036
rect 29112 30976 29176 30980
rect 29192 31036 29256 31040
rect 29192 30980 29196 31036
rect 29196 30980 29252 31036
rect 29252 30980 29256 31036
rect 29192 30976 29256 30980
rect 29272 31036 29336 31040
rect 29272 30980 29276 31036
rect 29276 30980 29332 31036
rect 29332 30980 29336 31036
rect 29272 30976 29336 30980
rect 29352 31036 29416 31040
rect 29352 30980 29356 31036
rect 29356 30980 29412 31036
rect 29412 30980 29416 31036
rect 29352 30976 29416 30980
rect 12216 30492 12280 30496
rect 12216 30436 12220 30492
rect 12220 30436 12276 30492
rect 12276 30436 12280 30492
rect 12216 30432 12280 30436
rect 12296 30492 12360 30496
rect 12296 30436 12300 30492
rect 12300 30436 12356 30492
rect 12356 30436 12360 30492
rect 12296 30432 12360 30436
rect 12376 30492 12440 30496
rect 12376 30436 12380 30492
rect 12380 30436 12436 30492
rect 12436 30436 12440 30492
rect 12376 30432 12440 30436
rect 12456 30492 12520 30496
rect 12456 30436 12460 30492
rect 12460 30436 12516 30492
rect 12516 30436 12520 30492
rect 12456 30432 12520 30436
rect 23480 30492 23544 30496
rect 23480 30436 23484 30492
rect 23484 30436 23540 30492
rect 23540 30436 23544 30492
rect 23480 30432 23544 30436
rect 23560 30492 23624 30496
rect 23560 30436 23564 30492
rect 23564 30436 23620 30492
rect 23620 30436 23624 30492
rect 23560 30432 23624 30436
rect 23640 30492 23704 30496
rect 23640 30436 23644 30492
rect 23644 30436 23700 30492
rect 23700 30436 23704 30492
rect 23640 30432 23704 30436
rect 23720 30492 23784 30496
rect 23720 30436 23724 30492
rect 23724 30436 23780 30492
rect 23780 30436 23784 30492
rect 23720 30432 23784 30436
rect 6584 29948 6648 29952
rect 6584 29892 6588 29948
rect 6588 29892 6644 29948
rect 6644 29892 6648 29948
rect 6584 29888 6648 29892
rect 6664 29948 6728 29952
rect 6664 29892 6668 29948
rect 6668 29892 6724 29948
rect 6724 29892 6728 29948
rect 6664 29888 6728 29892
rect 6744 29948 6808 29952
rect 6744 29892 6748 29948
rect 6748 29892 6804 29948
rect 6804 29892 6808 29948
rect 6744 29888 6808 29892
rect 6824 29948 6888 29952
rect 6824 29892 6828 29948
rect 6828 29892 6884 29948
rect 6884 29892 6888 29948
rect 6824 29888 6888 29892
rect 17848 29948 17912 29952
rect 17848 29892 17852 29948
rect 17852 29892 17908 29948
rect 17908 29892 17912 29948
rect 17848 29888 17912 29892
rect 17928 29948 17992 29952
rect 17928 29892 17932 29948
rect 17932 29892 17988 29948
rect 17988 29892 17992 29948
rect 17928 29888 17992 29892
rect 18008 29948 18072 29952
rect 18008 29892 18012 29948
rect 18012 29892 18068 29948
rect 18068 29892 18072 29948
rect 18008 29888 18072 29892
rect 18088 29948 18152 29952
rect 18088 29892 18092 29948
rect 18092 29892 18148 29948
rect 18148 29892 18152 29948
rect 18088 29888 18152 29892
rect 29112 29948 29176 29952
rect 29112 29892 29116 29948
rect 29116 29892 29172 29948
rect 29172 29892 29176 29948
rect 29112 29888 29176 29892
rect 29192 29948 29256 29952
rect 29192 29892 29196 29948
rect 29196 29892 29252 29948
rect 29252 29892 29256 29948
rect 29192 29888 29256 29892
rect 29272 29948 29336 29952
rect 29272 29892 29276 29948
rect 29276 29892 29332 29948
rect 29332 29892 29336 29948
rect 29272 29888 29336 29892
rect 29352 29948 29416 29952
rect 29352 29892 29356 29948
rect 29356 29892 29412 29948
rect 29412 29892 29416 29948
rect 29352 29888 29416 29892
rect 12216 29404 12280 29408
rect 12216 29348 12220 29404
rect 12220 29348 12276 29404
rect 12276 29348 12280 29404
rect 12216 29344 12280 29348
rect 12296 29404 12360 29408
rect 12296 29348 12300 29404
rect 12300 29348 12356 29404
rect 12356 29348 12360 29404
rect 12296 29344 12360 29348
rect 12376 29404 12440 29408
rect 12376 29348 12380 29404
rect 12380 29348 12436 29404
rect 12436 29348 12440 29404
rect 12376 29344 12440 29348
rect 12456 29404 12520 29408
rect 12456 29348 12460 29404
rect 12460 29348 12516 29404
rect 12516 29348 12520 29404
rect 12456 29344 12520 29348
rect 23480 29404 23544 29408
rect 23480 29348 23484 29404
rect 23484 29348 23540 29404
rect 23540 29348 23544 29404
rect 23480 29344 23544 29348
rect 23560 29404 23624 29408
rect 23560 29348 23564 29404
rect 23564 29348 23620 29404
rect 23620 29348 23624 29404
rect 23560 29344 23624 29348
rect 23640 29404 23704 29408
rect 23640 29348 23644 29404
rect 23644 29348 23700 29404
rect 23700 29348 23704 29404
rect 23640 29344 23704 29348
rect 23720 29404 23784 29408
rect 23720 29348 23724 29404
rect 23724 29348 23780 29404
rect 23780 29348 23784 29404
rect 23720 29344 23784 29348
rect 6584 28860 6648 28864
rect 6584 28804 6588 28860
rect 6588 28804 6644 28860
rect 6644 28804 6648 28860
rect 6584 28800 6648 28804
rect 6664 28860 6728 28864
rect 6664 28804 6668 28860
rect 6668 28804 6724 28860
rect 6724 28804 6728 28860
rect 6664 28800 6728 28804
rect 6744 28860 6808 28864
rect 6744 28804 6748 28860
rect 6748 28804 6804 28860
rect 6804 28804 6808 28860
rect 6744 28800 6808 28804
rect 6824 28860 6888 28864
rect 6824 28804 6828 28860
rect 6828 28804 6884 28860
rect 6884 28804 6888 28860
rect 6824 28800 6888 28804
rect 17848 28860 17912 28864
rect 17848 28804 17852 28860
rect 17852 28804 17908 28860
rect 17908 28804 17912 28860
rect 17848 28800 17912 28804
rect 17928 28860 17992 28864
rect 17928 28804 17932 28860
rect 17932 28804 17988 28860
rect 17988 28804 17992 28860
rect 17928 28800 17992 28804
rect 18008 28860 18072 28864
rect 18008 28804 18012 28860
rect 18012 28804 18068 28860
rect 18068 28804 18072 28860
rect 18008 28800 18072 28804
rect 18088 28860 18152 28864
rect 18088 28804 18092 28860
rect 18092 28804 18148 28860
rect 18148 28804 18152 28860
rect 18088 28800 18152 28804
rect 29112 28860 29176 28864
rect 29112 28804 29116 28860
rect 29116 28804 29172 28860
rect 29172 28804 29176 28860
rect 29112 28800 29176 28804
rect 29192 28860 29256 28864
rect 29192 28804 29196 28860
rect 29196 28804 29252 28860
rect 29252 28804 29256 28860
rect 29192 28800 29256 28804
rect 29272 28860 29336 28864
rect 29272 28804 29276 28860
rect 29276 28804 29332 28860
rect 29332 28804 29336 28860
rect 29272 28800 29336 28804
rect 29352 28860 29416 28864
rect 29352 28804 29356 28860
rect 29356 28804 29412 28860
rect 29412 28804 29416 28860
rect 29352 28800 29416 28804
rect 12216 28316 12280 28320
rect 12216 28260 12220 28316
rect 12220 28260 12276 28316
rect 12276 28260 12280 28316
rect 12216 28256 12280 28260
rect 12296 28316 12360 28320
rect 12296 28260 12300 28316
rect 12300 28260 12356 28316
rect 12356 28260 12360 28316
rect 12296 28256 12360 28260
rect 12376 28316 12440 28320
rect 12376 28260 12380 28316
rect 12380 28260 12436 28316
rect 12436 28260 12440 28316
rect 12376 28256 12440 28260
rect 12456 28316 12520 28320
rect 12456 28260 12460 28316
rect 12460 28260 12516 28316
rect 12516 28260 12520 28316
rect 12456 28256 12520 28260
rect 23480 28316 23544 28320
rect 23480 28260 23484 28316
rect 23484 28260 23540 28316
rect 23540 28260 23544 28316
rect 23480 28256 23544 28260
rect 23560 28316 23624 28320
rect 23560 28260 23564 28316
rect 23564 28260 23620 28316
rect 23620 28260 23624 28316
rect 23560 28256 23624 28260
rect 23640 28316 23704 28320
rect 23640 28260 23644 28316
rect 23644 28260 23700 28316
rect 23700 28260 23704 28316
rect 23640 28256 23704 28260
rect 23720 28316 23784 28320
rect 23720 28260 23724 28316
rect 23724 28260 23780 28316
rect 23780 28260 23784 28316
rect 23720 28256 23784 28260
rect 6584 27772 6648 27776
rect 6584 27716 6588 27772
rect 6588 27716 6644 27772
rect 6644 27716 6648 27772
rect 6584 27712 6648 27716
rect 6664 27772 6728 27776
rect 6664 27716 6668 27772
rect 6668 27716 6724 27772
rect 6724 27716 6728 27772
rect 6664 27712 6728 27716
rect 6744 27772 6808 27776
rect 6744 27716 6748 27772
rect 6748 27716 6804 27772
rect 6804 27716 6808 27772
rect 6744 27712 6808 27716
rect 6824 27772 6888 27776
rect 6824 27716 6828 27772
rect 6828 27716 6884 27772
rect 6884 27716 6888 27772
rect 6824 27712 6888 27716
rect 17848 27772 17912 27776
rect 17848 27716 17852 27772
rect 17852 27716 17908 27772
rect 17908 27716 17912 27772
rect 17848 27712 17912 27716
rect 17928 27772 17992 27776
rect 17928 27716 17932 27772
rect 17932 27716 17988 27772
rect 17988 27716 17992 27772
rect 17928 27712 17992 27716
rect 18008 27772 18072 27776
rect 18008 27716 18012 27772
rect 18012 27716 18068 27772
rect 18068 27716 18072 27772
rect 18008 27712 18072 27716
rect 18088 27772 18152 27776
rect 18088 27716 18092 27772
rect 18092 27716 18148 27772
rect 18148 27716 18152 27772
rect 18088 27712 18152 27716
rect 29112 27772 29176 27776
rect 29112 27716 29116 27772
rect 29116 27716 29172 27772
rect 29172 27716 29176 27772
rect 29112 27712 29176 27716
rect 29192 27772 29256 27776
rect 29192 27716 29196 27772
rect 29196 27716 29252 27772
rect 29252 27716 29256 27772
rect 29192 27712 29256 27716
rect 29272 27772 29336 27776
rect 29272 27716 29276 27772
rect 29276 27716 29332 27772
rect 29332 27716 29336 27772
rect 29272 27712 29336 27716
rect 29352 27772 29416 27776
rect 29352 27716 29356 27772
rect 29356 27716 29412 27772
rect 29412 27716 29416 27772
rect 29352 27712 29416 27716
rect 12216 27228 12280 27232
rect 12216 27172 12220 27228
rect 12220 27172 12276 27228
rect 12276 27172 12280 27228
rect 12216 27168 12280 27172
rect 12296 27228 12360 27232
rect 12296 27172 12300 27228
rect 12300 27172 12356 27228
rect 12356 27172 12360 27228
rect 12296 27168 12360 27172
rect 12376 27228 12440 27232
rect 12376 27172 12380 27228
rect 12380 27172 12436 27228
rect 12436 27172 12440 27228
rect 12376 27168 12440 27172
rect 12456 27228 12520 27232
rect 12456 27172 12460 27228
rect 12460 27172 12516 27228
rect 12516 27172 12520 27228
rect 12456 27168 12520 27172
rect 23480 27228 23544 27232
rect 23480 27172 23484 27228
rect 23484 27172 23540 27228
rect 23540 27172 23544 27228
rect 23480 27168 23544 27172
rect 23560 27228 23624 27232
rect 23560 27172 23564 27228
rect 23564 27172 23620 27228
rect 23620 27172 23624 27228
rect 23560 27168 23624 27172
rect 23640 27228 23704 27232
rect 23640 27172 23644 27228
rect 23644 27172 23700 27228
rect 23700 27172 23704 27228
rect 23640 27168 23704 27172
rect 23720 27228 23784 27232
rect 23720 27172 23724 27228
rect 23724 27172 23780 27228
rect 23780 27172 23784 27228
rect 23720 27168 23784 27172
rect 6584 26684 6648 26688
rect 6584 26628 6588 26684
rect 6588 26628 6644 26684
rect 6644 26628 6648 26684
rect 6584 26624 6648 26628
rect 6664 26684 6728 26688
rect 6664 26628 6668 26684
rect 6668 26628 6724 26684
rect 6724 26628 6728 26684
rect 6664 26624 6728 26628
rect 6744 26684 6808 26688
rect 6744 26628 6748 26684
rect 6748 26628 6804 26684
rect 6804 26628 6808 26684
rect 6744 26624 6808 26628
rect 6824 26684 6888 26688
rect 6824 26628 6828 26684
rect 6828 26628 6884 26684
rect 6884 26628 6888 26684
rect 6824 26624 6888 26628
rect 17848 26684 17912 26688
rect 17848 26628 17852 26684
rect 17852 26628 17908 26684
rect 17908 26628 17912 26684
rect 17848 26624 17912 26628
rect 17928 26684 17992 26688
rect 17928 26628 17932 26684
rect 17932 26628 17988 26684
rect 17988 26628 17992 26684
rect 17928 26624 17992 26628
rect 18008 26684 18072 26688
rect 18008 26628 18012 26684
rect 18012 26628 18068 26684
rect 18068 26628 18072 26684
rect 18008 26624 18072 26628
rect 18088 26684 18152 26688
rect 18088 26628 18092 26684
rect 18092 26628 18148 26684
rect 18148 26628 18152 26684
rect 18088 26624 18152 26628
rect 29112 26684 29176 26688
rect 29112 26628 29116 26684
rect 29116 26628 29172 26684
rect 29172 26628 29176 26684
rect 29112 26624 29176 26628
rect 29192 26684 29256 26688
rect 29192 26628 29196 26684
rect 29196 26628 29252 26684
rect 29252 26628 29256 26684
rect 29192 26624 29256 26628
rect 29272 26684 29336 26688
rect 29272 26628 29276 26684
rect 29276 26628 29332 26684
rect 29332 26628 29336 26684
rect 29272 26624 29336 26628
rect 29352 26684 29416 26688
rect 29352 26628 29356 26684
rect 29356 26628 29412 26684
rect 29412 26628 29416 26684
rect 29352 26624 29416 26628
rect 12216 26140 12280 26144
rect 12216 26084 12220 26140
rect 12220 26084 12276 26140
rect 12276 26084 12280 26140
rect 12216 26080 12280 26084
rect 12296 26140 12360 26144
rect 12296 26084 12300 26140
rect 12300 26084 12356 26140
rect 12356 26084 12360 26140
rect 12296 26080 12360 26084
rect 12376 26140 12440 26144
rect 12376 26084 12380 26140
rect 12380 26084 12436 26140
rect 12436 26084 12440 26140
rect 12376 26080 12440 26084
rect 12456 26140 12520 26144
rect 12456 26084 12460 26140
rect 12460 26084 12516 26140
rect 12516 26084 12520 26140
rect 12456 26080 12520 26084
rect 23480 26140 23544 26144
rect 23480 26084 23484 26140
rect 23484 26084 23540 26140
rect 23540 26084 23544 26140
rect 23480 26080 23544 26084
rect 23560 26140 23624 26144
rect 23560 26084 23564 26140
rect 23564 26084 23620 26140
rect 23620 26084 23624 26140
rect 23560 26080 23624 26084
rect 23640 26140 23704 26144
rect 23640 26084 23644 26140
rect 23644 26084 23700 26140
rect 23700 26084 23704 26140
rect 23640 26080 23704 26084
rect 23720 26140 23784 26144
rect 23720 26084 23724 26140
rect 23724 26084 23780 26140
rect 23780 26084 23784 26140
rect 23720 26080 23784 26084
rect 6584 25596 6648 25600
rect 6584 25540 6588 25596
rect 6588 25540 6644 25596
rect 6644 25540 6648 25596
rect 6584 25536 6648 25540
rect 6664 25596 6728 25600
rect 6664 25540 6668 25596
rect 6668 25540 6724 25596
rect 6724 25540 6728 25596
rect 6664 25536 6728 25540
rect 6744 25596 6808 25600
rect 6744 25540 6748 25596
rect 6748 25540 6804 25596
rect 6804 25540 6808 25596
rect 6744 25536 6808 25540
rect 6824 25596 6888 25600
rect 6824 25540 6828 25596
rect 6828 25540 6884 25596
rect 6884 25540 6888 25596
rect 6824 25536 6888 25540
rect 17848 25596 17912 25600
rect 17848 25540 17852 25596
rect 17852 25540 17908 25596
rect 17908 25540 17912 25596
rect 17848 25536 17912 25540
rect 17928 25596 17992 25600
rect 17928 25540 17932 25596
rect 17932 25540 17988 25596
rect 17988 25540 17992 25596
rect 17928 25536 17992 25540
rect 18008 25596 18072 25600
rect 18008 25540 18012 25596
rect 18012 25540 18068 25596
rect 18068 25540 18072 25596
rect 18008 25536 18072 25540
rect 18088 25596 18152 25600
rect 18088 25540 18092 25596
rect 18092 25540 18148 25596
rect 18148 25540 18152 25596
rect 18088 25536 18152 25540
rect 29112 25596 29176 25600
rect 29112 25540 29116 25596
rect 29116 25540 29172 25596
rect 29172 25540 29176 25596
rect 29112 25536 29176 25540
rect 29192 25596 29256 25600
rect 29192 25540 29196 25596
rect 29196 25540 29252 25596
rect 29252 25540 29256 25596
rect 29192 25536 29256 25540
rect 29272 25596 29336 25600
rect 29272 25540 29276 25596
rect 29276 25540 29332 25596
rect 29332 25540 29336 25596
rect 29272 25536 29336 25540
rect 29352 25596 29416 25600
rect 29352 25540 29356 25596
rect 29356 25540 29412 25596
rect 29412 25540 29416 25596
rect 29352 25536 29416 25540
rect 12216 25052 12280 25056
rect 12216 24996 12220 25052
rect 12220 24996 12276 25052
rect 12276 24996 12280 25052
rect 12216 24992 12280 24996
rect 12296 25052 12360 25056
rect 12296 24996 12300 25052
rect 12300 24996 12356 25052
rect 12356 24996 12360 25052
rect 12296 24992 12360 24996
rect 12376 25052 12440 25056
rect 12376 24996 12380 25052
rect 12380 24996 12436 25052
rect 12436 24996 12440 25052
rect 12376 24992 12440 24996
rect 12456 25052 12520 25056
rect 12456 24996 12460 25052
rect 12460 24996 12516 25052
rect 12516 24996 12520 25052
rect 12456 24992 12520 24996
rect 23480 25052 23544 25056
rect 23480 24996 23484 25052
rect 23484 24996 23540 25052
rect 23540 24996 23544 25052
rect 23480 24992 23544 24996
rect 23560 25052 23624 25056
rect 23560 24996 23564 25052
rect 23564 24996 23620 25052
rect 23620 24996 23624 25052
rect 23560 24992 23624 24996
rect 23640 25052 23704 25056
rect 23640 24996 23644 25052
rect 23644 24996 23700 25052
rect 23700 24996 23704 25052
rect 23640 24992 23704 24996
rect 23720 25052 23784 25056
rect 23720 24996 23724 25052
rect 23724 24996 23780 25052
rect 23780 24996 23784 25052
rect 23720 24992 23784 24996
rect 6584 24508 6648 24512
rect 6584 24452 6588 24508
rect 6588 24452 6644 24508
rect 6644 24452 6648 24508
rect 6584 24448 6648 24452
rect 6664 24508 6728 24512
rect 6664 24452 6668 24508
rect 6668 24452 6724 24508
rect 6724 24452 6728 24508
rect 6664 24448 6728 24452
rect 6744 24508 6808 24512
rect 6744 24452 6748 24508
rect 6748 24452 6804 24508
rect 6804 24452 6808 24508
rect 6744 24448 6808 24452
rect 6824 24508 6888 24512
rect 6824 24452 6828 24508
rect 6828 24452 6884 24508
rect 6884 24452 6888 24508
rect 6824 24448 6888 24452
rect 17848 24508 17912 24512
rect 17848 24452 17852 24508
rect 17852 24452 17908 24508
rect 17908 24452 17912 24508
rect 17848 24448 17912 24452
rect 17928 24508 17992 24512
rect 17928 24452 17932 24508
rect 17932 24452 17988 24508
rect 17988 24452 17992 24508
rect 17928 24448 17992 24452
rect 18008 24508 18072 24512
rect 18008 24452 18012 24508
rect 18012 24452 18068 24508
rect 18068 24452 18072 24508
rect 18008 24448 18072 24452
rect 18088 24508 18152 24512
rect 18088 24452 18092 24508
rect 18092 24452 18148 24508
rect 18148 24452 18152 24508
rect 18088 24448 18152 24452
rect 29112 24508 29176 24512
rect 29112 24452 29116 24508
rect 29116 24452 29172 24508
rect 29172 24452 29176 24508
rect 29112 24448 29176 24452
rect 29192 24508 29256 24512
rect 29192 24452 29196 24508
rect 29196 24452 29252 24508
rect 29252 24452 29256 24508
rect 29192 24448 29256 24452
rect 29272 24508 29336 24512
rect 29272 24452 29276 24508
rect 29276 24452 29332 24508
rect 29332 24452 29336 24508
rect 29272 24448 29336 24452
rect 29352 24508 29416 24512
rect 29352 24452 29356 24508
rect 29356 24452 29412 24508
rect 29412 24452 29416 24508
rect 29352 24448 29416 24452
rect 12216 23964 12280 23968
rect 12216 23908 12220 23964
rect 12220 23908 12276 23964
rect 12276 23908 12280 23964
rect 12216 23904 12280 23908
rect 12296 23964 12360 23968
rect 12296 23908 12300 23964
rect 12300 23908 12356 23964
rect 12356 23908 12360 23964
rect 12296 23904 12360 23908
rect 12376 23964 12440 23968
rect 12376 23908 12380 23964
rect 12380 23908 12436 23964
rect 12436 23908 12440 23964
rect 12376 23904 12440 23908
rect 12456 23964 12520 23968
rect 12456 23908 12460 23964
rect 12460 23908 12516 23964
rect 12516 23908 12520 23964
rect 12456 23904 12520 23908
rect 23480 23964 23544 23968
rect 23480 23908 23484 23964
rect 23484 23908 23540 23964
rect 23540 23908 23544 23964
rect 23480 23904 23544 23908
rect 23560 23964 23624 23968
rect 23560 23908 23564 23964
rect 23564 23908 23620 23964
rect 23620 23908 23624 23964
rect 23560 23904 23624 23908
rect 23640 23964 23704 23968
rect 23640 23908 23644 23964
rect 23644 23908 23700 23964
rect 23700 23908 23704 23964
rect 23640 23904 23704 23908
rect 23720 23964 23784 23968
rect 23720 23908 23724 23964
rect 23724 23908 23780 23964
rect 23780 23908 23784 23964
rect 23720 23904 23784 23908
rect 6584 23420 6648 23424
rect 6584 23364 6588 23420
rect 6588 23364 6644 23420
rect 6644 23364 6648 23420
rect 6584 23360 6648 23364
rect 6664 23420 6728 23424
rect 6664 23364 6668 23420
rect 6668 23364 6724 23420
rect 6724 23364 6728 23420
rect 6664 23360 6728 23364
rect 6744 23420 6808 23424
rect 6744 23364 6748 23420
rect 6748 23364 6804 23420
rect 6804 23364 6808 23420
rect 6744 23360 6808 23364
rect 6824 23420 6888 23424
rect 6824 23364 6828 23420
rect 6828 23364 6884 23420
rect 6884 23364 6888 23420
rect 6824 23360 6888 23364
rect 17848 23420 17912 23424
rect 17848 23364 17852 23420
rect 17852 23364 17908 23420
rect 17908 23364 17912 23420
rect 17848 23360 17912 23364
rect 17928 23420 17992 23424
rect 17928 23364 17932 23420
rect 17932 23364 17988 23420
rect 17988 23364 17992 23420
rect 17928 23360 17992 23364
rect 18008 23420 18072 23424
rect 18008 23364 18012 23420
rect 18012 23364 18068 23420
rect 18068 23364 18072 23420
rect 18008 23360 18072 23364
rect 18088 23420 18152 23424
rect 18088 23364 18092 23420
rect 18092 23364 18148 23420
rect 18148 23364 18152 23420
rect 18088 23360 18152 23364
rect 29112 23420 29176 23424
rect 29112 23364 29116 23420
rect 29116 23364 29172 23420
rect 29172 23364 29176 23420
rect 29112 23360 29176 23364
rect 29192 23420 29256 23424
rect 29192 23364 29196 23420
rect 29196 23364 29252 23420
rect 29252 23364 29256 23420
rect 29192 23360 29256 23364
rect 29272 23420 29336 23424
rect 29272 23364 29276 23420
rect 29276 23364 29332 23420
rect 29332 23364 29336 23420
rect 29272 23360 29336 23364
rect 29352 23420 29416 23424
rect 29352 23364 29356 23420
rect 29356 23364 29412 23420
rect 29412 23364 29416 23420
rect 29352 23360 29416 23364
rect 12216 22876 12280 22880
rect 12216 22820 12220 22876
rect 12220 22820 12276 22876
rect 12276 22820 12280 22876
rect 12216 22816 12280 22820
rect 12296 22876 12360 22880
rect 12296 22820 12300 22876
rect 12300 22820 12356 22876
rect 12356 22820 12360 22876
rect 12296 22816 12360 22820
rect 12376 22876 12440 22880
rect 12376 22820 12380 22876
rect 12380 22820 12436 22876
rect 12436 22820 12440 22876
rect 12376 22816 12440 22820
rect 12456 22876 12520 22880
rect 12456 22820 12460 22876
rect 12460 22820 12516 22876
rect 12516 22820 12520 22876
rect 12456 22816 12520 22820
rect 23480 22876 23544 22880
rect 23480 22820 23484 22876
rect 23484 22820 23540 22876
rect 23540 22820 23544 22876
rect 23480 22816 23544 22820
rect 23560 22876 23624 22880
rect 23560 22820 23564 22876
rect 23564 22820 23620 22876
rect 23620 22820 23624 22876
rect 23560 22816 23624 22820
rect 23640 22876 23704 22880
rect 23640 22820 23644 22876
rect 23644 22820 23700 22876
rect 23700 22820 23704 22876
rect 23640 22816 23704 22820
rect 23720 22876 23784 22880
rect 23720 22820 23724 22876
rect 23724 22820 23780 22876
rect 23780 22820 23784 22876
rect 23720 22816 23784 22820
rect 6584 22332 6648 22336
rect 6584 22276 6588 22332
rect 6588 22276 6644 22332
rect 6644 22276 6648 22332
rect 6584 22272 6648 22276
rect 6664 22332 6728 22336
rect 6664 22276 6668 22332
rect 6668 22276 6724 22332
rect 6724 22276 6728 22332
rect 6664 22272 6728 22276
rect 6744 22332 6808 22336
rect 6744 22276 6748 22332
rect 6748 22276 6804 22332
rect 6804 22276 6808 22332
rect 6744 22272 6808 22276
rect 6824 22332 6888 22336
rect 6824 22276 6828 22332
rect 6828 22276 6884 22332
rect 6884 22276 6888 22332
rect 6824 22272 6888 22276
rect 17848 22332 17912 22336
rect 17848 22276 17852 22332
rect 17852 22276 17908 22332
rect 17908 22276 17912 22332
rect 17848 22272 17912 22276
rect 17928 22332 17992 22336
rect 17928 22276 17932 22332
rect 17932 22276 17988 22332
rect 17988 22276 17992 22332
rect 17928 22272 17992 22276
rect 18008 22332 18072 22336
rect 18008 22276 18012 22332
rect 18012 22276 18068 22332
rect 18068 22276 18072 22332
rect 18008 22272 18072 22276
rect 18088 22332 18152 22336
rect 18088 22276 18092 22332
rect 18092 22276 18148 22332
rect 18148 22276 18152 22332
rect 18088 22272 18152 22276
rect 29112 22332 29176 22336
rect 29112 22276 29116 22332
rect 29116 22276 29172 22332
rect 29172 22276 29176 22332
rect 29112 22272 29176 22276
rect 29192 22332 29256 22336
rect 29192 22276 29196 22332
rect 29196 22276 29252 22332
rect 29252 22276 29256 22332
rect 29192 22272 29256 22276
rect 29272 22332 29336 22336
rect 29272 22276 29276 22332
rect 29276 22276 29332 22332
rect 29332 22276 29336 22332
rect 29272 22272 29336 22276
rect 29352 22332 29416 22336
rect 29352 22276 29356 22332
rect 29356 22276 29412 22332
rect 29412 22276 29416 22332
rect 29352 22272 29416 22276
rect 12216 21788 12280 21792
rect 12216 21732 12220 21788
rect 12220 21732 12276 21788
rect 12276 21732 12280 21788
rect 12216 21728 12280 21732
rect 12296 21788 12360 21792
rect 12296 21732 12300 21788
rect 12300 21732 12356 21788
rect 12356 21732 12360 21788
rect 12296 21728 12360 21732
rect 12376 21788 12440 21792
rect 12376 21732 12380 21788
rect 12380 21732 12436 21788
rect 12436 21732 12440 21788
rect 12376 21728 12440 21732
rect 12456 21788 12520 21792
rect 12456 21732 12460 21788
rect 12460 21732 12516 21788
rect 12516 21732 12520 21788
rect 12456 21728 12520 21732
rect 23480 21788 23544 21792
rect 23480 21732 23484 21788
rect 23484 21732 23540 21788
rect 23540 21732 23544 21788
rect 23480 21728 23544 21732
rect 23560 21788 23624 21792
rect 23560 21732 23564 21788
rect 23564 21732 23620 21788
rect 23620 21732 23624 21788
rect 23560 21728 23624 21732
rect 23640 21788 23704 21792
rect 23640 21732 23644 21788
rect 23644 21732 23700 21788
rect 23700 21732 23704 21788
rect 23640 21728 23704 21732
rect 23720 21788 23784 21792
rect 23720 21732 23724 21788
rect 23724 21732 23780 21788
rect 23780 21732 23784 21788
rect 23720 21728 23784 21732
rect 6584 21244 6648 21248
rect 6584 21188 6588 21244
rect 6588 21188 6644 21244
rect 6644 21188 6648 21244
rect 6584 21184 6648 21188
rect 6664 21244 6728 21248
rect 6664 21188 6668 21244
rect 6668 21188 6724 21244
rect 6724 21188 6728 21244
rect 6664 21184 6728 21188
rect 6744 21244 6808 21248
rect 6744 21188 6748 21244
rect 6748 21188 6804 21244
rect 6804 21188 6808 21244
rect 6744 21184 6808 21188
rect 6824 21244 6888 21248
rect 6824 21188 6828 21244
rect 6828 21188 6884 21244
rect 6884 21188 6888 21244
rect 6824 21184 6888 21188
rect 17848 21244 17912 21248
rect 17848 21188 17852 21244
rect 17852 21188 17908 21244
rect 17908 21188 17912 21244
rect 17848 21184 17912 21188
rect 17928 21244 17992 21248
rect 17928 21188 17932 21244
rect 17932 21188 17988 21244
rect 17988 21188 17992 21244
rect 17928 21184 17992 21188
rect 18008 21244 18072 21248
rect 18008 21188 18012 21244
rect 18012 21188 18068 21244
rect 18068 21188 18072 21244
rect 18008 21184 18072 21188
rect 18088 21244 18152 21248
rect 18088 21188 18092 21244
rect 18092 21188 18148 21244
rect 18148 21188 18152 21244
rect 18088 21184 18152 21188
rect 29112 21244 29176 21248
rect 29112 21188 29116 21244
rect 29116 21188 29172 21244
rect 29172 21188 29176 21244
rect 29112 21184 29176 21188
rect 29192 21244 29256 21248
rect 29192 21188 29196 21244
rect 29196 21188 29252 21244
rect 29252 21188 29256 21244
rect 29192 21184 29256 21188
rect 29272 21244 29336 21248
rect 29272 21188 29276 21244
rect 29276 21188 29332 21244
rect 29332 21188 29336 21244
rect 29272 21184 29336 21188
rect 29352 21244 29416 21248
rect 29352 21188 29356 21244
rect 29356 21188 29412 21244
rect 29412 21188 29416 21244
rect 29352 21184 29416 21188
rect 12216 20700 12280 20704
rect 12216 20644 12220 20700
rect 12220 20644 12276 20700
rect 12276 20644 12280 20700
rect 12216 20640 12280 20644
rect 12296 20700 12360 20704
rect 12296 20644 12300 20700
rect 12300 20644 12356 20700
rect 12356 20644 12360 20700
rect 12296 20640 12360 20644
rect 12376 20700 12440 20704
rect 12376 20644 12380 20700
rect 12380 20644 12436 20700
rect 12436 20644 12440 20700
rect 12376 20640 12440 20644
rect 12456 20700 12520 20704
rect 12456 20644 12460 20700
rect 12460 20644 12516 20700
rect 12516 20644 12520 20700
rect 12456 20640 12520 20644
rect 23480 20700 23544 20704
rect 23480 20644 23484 20700
rect 23484 20644 23540 20700
rect 23540 20644 23544 20700
rect 23480 20640 23544 20644
rect 23560 20700 23624 20704
rect 23560 20644 23564 20700
rect 23564 20644 23620 20700
rect 23620 20644 23624 20700
rect 23560 20640 23624 20644
rect 23640 20700 23704 20704
rect 23640 20644 23644 20700
rect 23644 20644 23700 20700
rect 23700 20644 23704 20700
rect 23640 20640 23704 20644
rect 23720 20700 23784 20704
rect 23720 20644 23724 20700
rect 23724 20644 23780 20700
rect 23780 20644 23784 20700
rect 23720 20640 23784 20644
rect 6584 20156 6648 20160
rect 6584 20100 6588 20156
rect 6588 20100 6644 20156
rect 6644 20100 6648 20156
rect 6584 20096 6648 20100
rect 6664 20156 6728 20160
rect 6664 20100 6668 20156
rect 6668 20100 6724 20156
rect 6724 20100 6728 20156
rect 6664 20096 6728 20100
rect 6744 20156 6808 20160
rect 6744 20100 6748 20156
rect 6748 20100 6804 20156
rect 6804 20100 6808 20156
rect 6744 20096 6808 20100
rect 6824 20156 6888 20160
rect 6824 20100 6828 20156
rect 6828 20100 6884 20156
rect 6884 20100 6888 20156
rect 6824 20096 6888 20100
rect 17848 20156 17912 20160
rect 17848 20100 17852 20156
rect 17852 20100 17908 20156
rect 17908 20100 17912 20156
rect 17848 20096 17912 20100
rect 17928 20156 17992 20160
rect 17928 20100 17932 20156
rect 17932 20100 17988 20156
rect 17988 20100 17992 20156
rect 17928 20096 17992 20100
rect 18008 20156 18072 20160
rect 18008 20100 18012 20156
rect 18012 20100 18068 20156
rect 18068 20100 18072 20156
rect 18008 20096 18072 20100
rect 18088 20156 18152 20160
rect 18088 20100 18092 20156
rect 18092 20100 18148 20156
rect 18148 20100 18152 20156
rect 18088 20096 18152 20100
rect 29112 20156 29176 20160
rect 29112 20100 29116 20156
rect 29116 20100 29172 20156
rect 29172 20100 29176 20156
rect 29112 20096 29176 20100
rect 29192 20156 29256 20160
rect 29192 20100 29196 20156
rect 29196 20100 29252 20156
rect 29252 20100 29256 20156
rect 29192 20096 29256 20100
rect 29272 20156 29336 20160
rect 29272 20100 29276 20156
rect 29276 20100 29332 20156
rect 29332 20100 29336 20156
rect 29272 20096 29336 20100
rect 29352 20156 29416 20160
rect 29352 20100 29356 20156
rect 29356 20100 29412 20156
rect 29412 20100 29416 20156
rect 29352 20096 29416 20100
rect 12216 19612 12280 19616
rect 12216 19556 12220 19612
rect 12220 19556 12276 19612
rect 12276 19556 12280 19612
rect 12216 19552 12280 19556
rect 12296 19612 12360 19616
rect 12296 19556 12300 19612
rect 12300 19556 12356 19612
rect 12356 19556 12360 19612
rect 12296 19552 12360 19556
rect 12376 19612 12440 19616
rect 12376 19556 12380 19612
rect 12380 19556 12436 19612
rect 12436 19556 12440 19612
rect 12376 19552 12440 19556
rect 12456 19612 12520 19616
rect 12456 19556 12460 19612
rect 12460 19556 12516 19612
rect 12516 19556 12520 19612
rect 12456 19552 12520 19556
rect 23480 19612 23544 19616
rect 23480 19556 23484 19612
rect 23484 19556 23540 19612
rect 23540 19556 23544 19612
rect 23480 19552 23544 19556
rect 23560 19612 23624 19616
rect 23560 19556 23564 19612
rect 23564 19556 23620 19612
rect 23620 19556 23624 19612
rect 23560 19552 23624 19556
rect 23640 19612 23704 19616
rect 23640 19556 23644 19612
rect 23644 19556 23700 19612
rect 23700 19556 23704 19612
rect 23640 19552 23704 19556
rect 23720 19612 23784 19616
rect 23720 19556 23724 19612
rect 23724 19556 23780 19612
rect 23780 19556 23784 19612
rect 23720 19552 23784 19556
rect 6584 19068 6648 19072
rect 6584 19012 6588 19068
rect 6588 19012 6644 19068
rect 6644 19012 6648 19068
rect 6584 19008 6648 19012
rect 6664 19068 6728 19072
rect 6664 19012 6668 19068
rect 6668 19012 6724 19068
rect 6724 19012 6728 19068
rect 6664 19008 6728 19012
rect 6744 19068 6808 19072
rect 6744 19012 6748 19068
rect 6748 19012 6804 19068
rect 6804 19012 6808 19068
rect 6744 19008 6808 19012
rect 6824 19068 6888 19072
rect 6824 19012 6828 19068
rect 6828 19012 6884 19068
rect 6884 19012 6888 19068
rect 6824 19008 6888 19012
rect 17848 19068 17912 19072
rect 17848 19012 17852 19068
rect 17852 19012 17908 19068
rect 17908 19012 17912 19068
rect 17848 19008 17912 19012
rect 17928 19068 17992 19072
rect 17928 19012 17932 19068
rect 17932 19012 17988 19068
rect 17988 19012 17992 19068
rect 17928 19008 17992 19012
rect 18008 19068 18072 19072
rect 18008 19012 18012 19068
rect 18012 19012 18068 19068
rect 18068 19012 18072 19068
rect 18008 19008 18072 19012
rect 18088 19068 18152 19072
rect 18088 19012 18092 19068
rect 18092 19012 18148 19068
rect 18148 19012 18152 19068
rect 18088 19008 18152 19012
rect 29112 19068 29176 19072
rect 29112 19012 29116 19068
rect 29116 19012 29172 19068
rect 29172 19012 29176 19068
rect 29112 19008 29176 19012
rect 29192 19068 29256 19072
rect 29192 19012 29196 19068
rect 29196 19012 29252 19068
rect 29252 19012 29256 19068
rect 29192 19008 29256 19012
rect 29272 19068 29336 19072
rect 29272 19012 29276 19068
rect 29276 19012 29332 19068
rect 29332 19012 29336 19068
rect 29272 19008 29336 19012
rect 29352 19068 29416 19072
rect 29352 19012 29356 19068
rect 29356 19012 29412 19068
rect 29412 19012 29416 19068
rect 29352 19008 29416 19012
rect 12216 18524 12280 18528
rect 12216 18468 12220 18524
rect 12220 18468 12276 18524
rect 12276 18468 12280 18524
rect 12216 18464 12280 18468
rect 12296 18524 12360 18528
rect 12296 18468 12300 18524
rect 12300 18468 12356 18524
rect 12356 18468 12360 18524
rect 12296 18464 12360 18468
rect 12376 18524 12440 18528
rect 12376 18468 12380 18524
rect 12380 18468 12436 18524
rect 12436 18468 12440 18524
rect 12376 18464 12440 18468
rect 12456 18524 12520 18528
rect 12456 18468 12460 18524
rect 12460 18468 12516 18524
rect 12516 18468 12520 18524
rect 12456 18464 12520 18468
rect 23480 18524 23544 18528
rect 23480 18468 23484 18524
rect 23484 18468 23540 18524
rect 23540 18468 23544 18524
rect 23480 18464 23544 18468
rect 23560 18524 23624 18528
rect 23560 18468 23564 18524
rect 23564 18468 23620 18524
rect 23620 18468 23624 18524
rect 23560 18464 23624 18468
rect 23640 18524 23704 18528
rect 23640 18468 23644 18524
rect 23644 18468 23700 18524
rect 23700 18468 23704 18524
rect 23640 18464 23704 18468
rect 23720 18524 23784 18528
rect 23720 18468 23724 18524
rect 23724 18468 23780 18524
rect 23780 18468 23784 18524
rect 23720 18464 23784 18468
rect 6584 17980 6648 17984
rect 6584 17924 6588 17980
rect 6588 17924 6644 17980
rect 6644 17924 6648 17980
rect 6584 17920 6648 17924
rect 6664 17980 6728 17984
rect 6664 17924 6668 17980
rect 6668 17924 6724 17980
rect 6724 17924 6728 17980
rect 6664 17920 6728 17924
rect 6744 17980 6808 17984
rect 6744 17924 6748 17980
rect 6748 17924 6804 17980
rect 6804 17924 6808 17980
rect 6744 17920 6808 17924
rect 6824 17980 6888 17984
rect 6824 17924 6828 17980
rect 6828 17924 6884 17980
rect 6884 17924 6888 17980
rect 6824 17920 6888 17924
rect 17848 17980 17912 17984
rect 17848 17924 17852 17980
rect 17852 17924 17908 17980
rect 17908 17924 17912 17980
rect 17848 17920 17912 17924
rect 17928 17980 17992 17984
rect 17928 17924 17932 17980
rect 17932 17924 17988 17980
rect 17988 17924 17992 17980
rect 17928 17920 17992 17924
rect 18008 17980 18072 17984
rect 18008 17924 18012 17980
rect 18012 17924 18068 17980
rect 18068 17924 18072 17980
rect 18008 17920 18072 17924
rect 18088 17980 18152 17984
rect 18088 17924 18092 17980
rect 18092 17924 18148 17980
rect 18148 17924 18152 17980
rect 18088 17920 18152 17924
rect 29112 17980 29176 17984
rect 29112 17924 29116 17980
rect 29116 17924 29172 17980
rect 29172 17924 29176 17980
rect 29112 17920 29176 17924
rect 29192 17980 29256 17984
rect 29192 17924 29196 17980
rect 29196 17924 29252 17980
rect 29252 17924 29256 17980
rect 29192 17920 29256 17924
rect 29272 17980 29336 17984
rect 29272 17924 29276 17980
rect 29276 17924 29332 17980
rect 29332 17924 29336 17980
rect 29272 17920 29336 17924
rect 29352 17980 29416 17984
rect 29352 17924 29356 17980
rect 29356 17924 29412 17980
rect 29412 17924 29416 17980
rect 29352 17920 29416 17924
rect 12216 17436 12280 17440
rect 12216 17380 12220 17436
rect 12220 17380 12276 17436
rect 12276 17380 12280 17436
rect 12216 17376 12280 17380
rect 12296 17436 12360 17440
rect 12296 17380 12300 17436
rect 12300 17380 12356 17436
rect 12356 17380 12360 17436
rect 12296 17376 12360 17380
rect 12376 17436 12440 17440
rect 12376 17380 12380 17436
rect 12380 17380 12436 17436
rect 12436 17380 12440 17436
rect 12376 17376 12440 17380
rect 12456 17436 12520 17440
rect 12456 17380 12460 17436
rect 12460 17380 12516 17436
rect 12516 17380 12520 17436
rect 12456 17376 12520 17380
rect 23480 17436 23544 17440
rect 23480 17380 23484 17436
rect 23484 17380 23540 17436
rect 23540 17380 23544 17436
rect 23480 17376 23544 17380
rect 23560 17436 23624 17440
rect 23560 17380 23564 17436
rect 23564 17380 23620 17436
rect 23620 17380 23624 17436
rect 23560 17376 23624 17380
rect 23640 17436 23704 17440
rect 23640 17380 23644 17436
rect 23644 17380 23700 17436
rect 23700 17380 23704 17436
rect 23640 17376 23704 17380
rect 23720 17436 23784 17440
rect 23720 17380 23724 17436
rect 23724 17380 23780 17436
rect 23780 17380 23784 17436
rect 23720 17376 23784 17380
rect 6584 16892 6648 16896
rect 6584 16836 6588 16892
rect 6588 16836 6644 16892
rect 6644 16836 6648 16892
rect 6584 16832 6648 16836
rect 6664 16892 6728 16896
rect 6664 16836 6668 16892
rect 6668 16836 6724 16892
rect 6724 16836 6728 16892
rect 6664 16832 6728 16836
rect 6744 16892 6808 16896
rect 6744 16836 6748 16892
rect 6748 16836 6804 16892
rect 6804 16836 6808 16892
rect 6744 16832 6808 16836
rect 6824 16892 6888 16896
rect 6824 16836 6828 16892
rect 6828 16836 6884 16892
rect 6884 16836 6888 16892
rect 6824 16832 6888 16836
rect 17848 16892 17912 16896
rect 17848 16836 17852 16892
rect 17852 16836 17908 16892
rect 17908 16836 17912 16892
rect 17848 16832 17912 16836
rect 17928 16892 17992 16896
rect 17928 16836 17932 16892
rect 17932 16836 17988 16892
rect 17988 16836 17992 16892
rect 17928 16832 17992 16836
rect 18008 16892 18072 16896
rect 18008 16836 18012 16892
rect 18012 16836 18068 16892
rect 18068 16836 18072 16892
rect 18008 16832 18072 16836
rect 18088 16892 18152 16896
rect 18088 16836 18092 16892
rect 18092 16836 18148 16892
rect 18148 16836 18152 16892
rect 18088 16832 18152 16836
rect 29112 16892 29176 16896
rect 29112 16836 29116 16892
rect 29116 16836 29172 16892
rect 29172 16836 29176 16892
rect 29112 16832 29176 16836
rect 29192 16892 29256 16896
rect 29192 16836 29196 16892
rect 29196 16836 29252 16892
rect 29252 16836 29256 16892
rect 29192 16832 29256 16836
rect 29272 16892 29336 16896
rect 29272 16836 29276 16892
rect 29276 16836 29332 16892
rect 29332 16836 29336 16892
rect 29272 16832 29336 16836
rect 29352 16892 29416 16896
rect 29352 16836 29356 16892
rect 29356 16836 29412 16892
rect 29412 16836 29416 16892
rect 29352 16832 29416 16836
rect 12216 16348 12280 16352
rect 12216 16292 12220 16348
rect 12220 16292 12276 16348
rect 12276 16292 12280 16348
rect 12216 16288 12280 16292
rect 12296 16348 12360 16352
rect 12296 16292 12300 16348
rect 12300 16292 12356 16348
rect 12356 16292 12360 16348
rect 12296 16288 12360 16292
rect 12376 16348 12440 16352
rect 12376 16292 12380 16348
rect 12380 16292 12436 16348
rect 12436 16292 12440 16348
rect 12376 16288 12440 16292
rect 12456 16348 12520 16352
rect 12456 16292 12460 16348
rect 12460 16292 12516 16348
rect 12516 16292 12520 16348
rect 12456 16288 12520 16292
rect 23480 16348 23544 16352
rect 23480 16292 23484 16348
rect 23484 16292 23540 16348
rect 23540 16292 23544 16348
rect 23480 16288 23544 16292
rect 23560 16348 23624 16352
rect 23560 16292 23564 16348
rect 23564 16292 23620 16348
rect 23620 16292 23624 16348
rect 23560 16288 23624 16292
rect 23640 16348 23704 16352
rect 23640 16292 23644 16348
rect 23644 16292 23700 16348
rect 23700 16292 23704 16348
rect 23640 16288 23704 16292
rect 23720 16348 23784 16352
rect 23720 16292 23724 16348
rect 23724 16292 23780 16348
rect 23780 16292 23784 16348
rect 23720 16288 23784 16292
rect 6584 15804 6648 15808
rect 6584 15748 6588 15804
rect 6588 15748 6644 15804
rect 6644 15748 6648 15804
rect 6584 15744 6648 15748
rect 6664 15804 6728 15808
rect 6664 15748 6668 15804
rect 6668 15748 6724 15804
rect 6724 15748 6728 15804
rect 6664 15744 6728 15748
rect 6744 15804 6808 15808
rect 6744 15748 6748 15804
rect 6748 15748 6804 15804
rect 6804 15748 6808 15804
rect 6744 15744 6808 15748
rect 6824 15804 6888 15808
rect 6824 15748 6828 15804
rect 6828 15748 6884 15804
rect 6884 15748 6888 15804
rect 6824 15744 6888 15748
rect 17848 15804 17912 15808
rect 17848 15748 17852 15804
rect 17852 15748 17908 15804
rect 17908 15748 17912 15804
rect 17848 15744 17912 15748
rect 17928 15804 17992 15808
rect 17928 15748 17932 15804
rect 17932 15748 17988 15804
rect 17988 15748 17992 15804
rect 17928 15744 17992 15748
rect 18008 15804 18072 15808
rect 18008 15748 18012 15804
rect 18012 15748 18068 15804
rect 18068 15748 18072 15804
rect 18008 15744 18072 15748
rect 18088 15804 18152 15808
rect 18088 15748 18092 15804
rect 18092 15748 18148 15804
rect 18148 15748 18152 15804
rect 18088 15744 18152 15748
rect 29112 15804 29176 15808
rect 29112 15748 29116 15804
rect 29116 15748 29172 15804
rect 29172 15748 29176 15804
rect 29112 15744 29176 15748
rect 29192 15804 29256 15808
rect 29192 15748 29196 15804
rect 29196 15748 29252 15804
rect 29252 15748 29256 15804
rect 29192 15744 29256 15748
rect 29272 15804 29336 15808
rect 29272 15748 29276 15804
rect 29276 15748 29332 15804
rect 29332 15748 29336 15804
rect 29272 15744 29336 15748
rect 29352 15804 29416 15808
rect 29352 15748 29356 15804
rect 29356 15748 29412 15804
rect 29412 15748 29416 15804
rect 29352 15744 29416 15748
rect 12216 15260 12280 15264
rect 12216 15204 12220 15260
rect 12220 15204 12276 15260
rect 12276 15204 12280 15260
rect 12216 15200 12280 15204
rect 12296 15260 12360 15264
rect 12296 15204 12300 15260
rect 12300 15204 12356 15260
rect 12356 15204 12360 15260
rect 12296 15200 12360 15204
rect 12376 15260 12440 15264
rect 12376 15204 12380 15260
rect 12380 15204 12436 15260
rect 12436 15204 12440 15260
rect 12376 15200 12440 15204
rect 12456 15260 12520 15264
rect 12456 15204 12460 15260
rect 12460 15204 12516 15260
rect 12516 15204 12520 15260
rect 12456 15200 12520 15204
rect 23480 15260 23544 15264
rect 23480 15204 23484 15260
rect 23484 15204 23540 15260
rect 23540 15204 23544 15260
rect 23480 15200 23544 15204
rect 23560 15260 23624 15264
rect 23560 15204 23564 15260
rect 23564 15204 23620 15260
rect 23620 15204 23624 15260
rect 23560 15200 23624 15204
rect 23640 15260 23704 15264
rect 23640 15204 23644 15260
rect 23644 15204 23700 15260
rect 23700 15204 23704 15260
rect 23640 15200 23704 15204
rect 23720 15260 23784 15264
rect 23720 15204 23724 15260
rect 23724 15204 23780 15260
rect 23780 15204 23784 15260
rect 23720 15200 23784 15204
rect 6584 14716 6648 14720
rect 6584 14660 6588 14716
rect 6588 14660 6644 14716
rect 6644 14660 6648 14716
rect 6584 14656 6648 14660
rect 6664 14716 6728 14720
rect 6664 14660 6668 14716
rect 6668 14660 6724 14716
rect 6724 14660 6728 14716
rect 6664 14656 6728 14660
rect 6744 14716 6808 14720
rect 6744 14660 6748 14716
rect 6748 14660 6804 14716
rect 6804 14660 6808 14716
rect 6744 14656 6808 14660
rect 6824 14716 6888 14720
rect 6824 14660 6828 14716
rect 6828 14660 6884 14716
rect 6884 14660 6888 14716
rect 6824 14656 6888 14660
rect 17848 14716 17912 14720
rect 17848 14660 17852 14716
rect 17852 14660 17908 14716
rect 17908 14660 17912 14716
rect 17848 14656 17912 14660
rect 17928 14716 17992 14720
rect 17928 14660 17932 14716
rect 17932 14660 17988 14716
rect 17988 14660 17992 14716
rect 17928 14656 17992 14660
rect 18008 14716 18072 14720
rect 18008 14660 18012 14716
rect 18012 14660 18068 14716
rect 18068 14660 18072 14716
rect 18008 14656 18072 14660
rect 18088 14716 18152 14720
rect 18088 14660 18092 14716
rect 18092 14660 18148 14716
rect 18148 14660 18152 14716
rect 18088 14656 18152 14660
rect 29112 14716 29176 14720
rect 29112 14660 29116 14716
rect 29116 14660 29172 14716
rect 29172 14660 29176 14716
rect 29112 14656 29176 14660
rect 29192 14716 29256 14720
rect 29192 14660 29196 14716
rect 29196 14660 29252 14716
rect 29252 14660 29256 14716
rect 29192 14656 29256 14660
rect 29272 14716 29336 14720
rect 29272 14660 29276 14716
rect 29276 14660 29332 14716
rect 29332 14660 29336 14716
rect 29272 14656 29336 14660
rect 29352 14716 29416 14720
rect 29352 14660 29356 14716
rect 29356 14660 29412 14716
rect 29412 14660 29416 14716
rect 29352 14656 29416 14660
rect 12216 14172 12280 14176
rect 12216 14116 12220 14172
rect 12220 14116 12276 14172
rect 12276 14116 12280 14172
rect 12216 14112 12280 14116
rect 12296 14172 12360 14176
rect 12296 14116 12300 14172
rect 12300 14116 12356 14172
rect 12356 14116 12360 14172
rect 12296 14112 12360 14116
rect 12376 14172 12440 14176
rect 12376 14116 12380 14172
rect 12380 14116 12436 14172
rect 12436 14116 12440 14172
rect 12376 14112 12440 14116
rect 12456 14172 12520 14176
rect 12456 14116 12460 14172
rect 12460 14116 12516 14172
rect 12516 14116 12520 14172
rect 12456 14112 12520 14116
rect 23480 14172 23544 14176
rect 23480 14116 23484 14172
rect 23484 14116 23540 14172
rect 23540 14116 23544 14172
rect 23480 14112 23544 14116
rect 23560 14172 23624 14176
rect 23560 14116 23564 14172
rect 23564 14116 23620 14172
rect 23620 14116 23624 14172
rect 23560 14112 23624 14116
rect 23640 14172 23704 14176
rect 23640 14116 23644 14172
rect 23644 14116 23700 14172
rect 23700 14116 23704 14172
rect 23640 14112 23704 14116
rect 23720 14172 23784 14176
rect 23720 14116 23724 14172
rect 23724 14116 23780 14172
rect 23780 14116 23784 14172
rect 23720 14112 23784 14116
rect 6584 13628 6648 13632
rect 6584 13572 6588 13628
rect 6588 13572 6644 13628
rect 6644 13572 6648 13628
rect 6584 13568 6648 13572
rect 6664 13628 6728 13632
rect 6664 13572 6668 13628
rect 6668 13572 6724 13628
rect 6724 13572 6728 13628
rect 6664 13568 6728 13572
rect 6744 13628 6808 13632
rect 6744 13572 6748 13628
rect 6748 13572 6804 13628
rect 6804 13572 6808 13628
rect 6744 13568 6808 13572
rect 6824 13628 6888 13632
rect 6824 13572 6828 13628
rect 6828 13572 6884 13628
rect 6884 13572 6888 13628
rect 6824 13568 6888 13572
rect 17848 13628 17912 13632
rect 17848 13572 17852 13628
rect 17852 13572 17908 13628
rect 17908 13572 17912 13628
rect 17848 13568 17912 13572
rect 17928 13628 17992 13632
rect 17928 13572 17932 13628
rect 17932 13572 17988 13628
rect 17988 13572 17992 13628
rect 17928 13568 17992 13572
rect 18008 13628 18072 13632
rect 18008 13572 18012 13628
rect 18012 13572 18068 13628
rect 18068 13572 18072 13628
rect 18008 13568 18072 13572
rect 18088 13628 18152 13632
rect 18088 13572 18092 13628
rect 18092 13572 18148 13628
rect 18148 13572 18152 13628
rect 18088 13568 18152 13572
rect 29112 13628 29176 13632
rect 29112 13572 29116 13628
rect 29116 13572 29172 13628
rect 29172 13572 29176 13628
rect 29112 13568 29176 13572
rect 29192 13628 29256 13632
rect 29192 13572 29196 13628
rect 29196 13572 29252 13628
rect 29252 13572 29256 13628
rect 29192 13568 29256 13572
rect 29272 13628 29336 13632
rect 29272 13572 29276 13628
rect 29276 13572 29332 13628
rect 29332 13572 29336 13628
rect 29272 13568 29336 13572
rect 29352 13628 29416 13632
rect 29352 13572 29356 13628
rect 29356 13572 29412 13628
rect 29412 13572 29416 13628
rect 29352 13568 29416 13572
rect 12216 13084 12280 13088
rect 12216 13028 12220 13084
rect 12220 13028 12276 13084
rect 12276 13028 12280 13084
rect 12216 13024 12280 13028
rect 12296 13084 12360 13088
rect 12296 13028 12300 13084
rect 12300 13028 12356 13084
rect 12356 13028 12360 13084
rect 12296 13024 12360 13028
rect 12376 13084 12440 13088
rect 12376 13028 12380 13084
rect 12380 13028 12436 13084
rect 12436 13028 12440 13084
rect 12376 13024 12440 13028
rect 12456 13084 12520 13088
rect 12456 13028 12460 13084
rect 12460 13028 12516 13084
rect 12516 13028 12520 13084
rect 12456 13024 12520 13028
rect 23480 13084 23544 13088
rect 23480 13028 23484 13084
rect 23484 13028 23540 13084
rect 23540 13028 23544 13084
rect 23480 13024 23544 13028
rect 23560 13084 23624 13088
rect 23560 13028 23564 13084
rect 23564 13028 23620 13084
rect 23620 13028 23624 13084
rect 23560 13024 23624 13028
rect 23640 13084 23704 13088
rect 23640 13028 23644 13084
rect 23644 13028 23700 13084
rect 23700 13028 23704 13084
rect 23640 13024 23704 13028
rect 23720 13084 23784 13088
rect 23720 13028 23724 13084
rect 23724 13028 23780 13084
rect 23780 13028 23784 13084
rect 23720 13024 23784 13028
rect 6584 12540 6648 12544
rect 6584 12484 6588 12540
rect 6588 12484 6644 12540
rect 6644 12484 6648 12540
rect 6584 12480 6648 12484
rect 6664 12540 6728 12544
rect 6664 12484 6668 12540
rect 6668 12484 6724 12540
rect 6724 12484 6728 12540
rect 6664 12480 6728 12484
rect 6744 12540 6808 12544
rect 6744 12484 6748 12540
rect 6748 12484 6804 12540
rect 6804 12484 6808 12540
rect 6744 12480 6808 12484
rect 6824 12540 6888 12544
rect 6824 12484 6828 12540
rect 6828 12484 6884 12540
rect 6884 12484 6888 12540
rect 6824 12480 6888 12484
rect 17848 12540 17912 12544
rect 17848 12484 17852 12540
rect 17852 12484 17908 12540
rect 17908 12484 17912 12540
rect 17848 12480 17912 12484
rect 17928 12540 17992 12544
rect 17928 12484 17932 12540
rect 17932 12484 17988 12540
rect 17988 12484 17992 12540
rect 17928 12480 17992 12484
rect 18008 12540 18072 12544
rect 18008 12484 18012 12540
rect 18012 12484 18068 12540
rect 18068 12484 18072 12540
rect 18008 12480 18072 12484
rect 18088 12540 18152 12544
rect 18088 12484 18092 12540
rect 18092 12484 18148 12540
rect 18148 12484 18152 12540
rect 18088 12480 18152 12484
rect 29112 12540 29176 12544
rect 29112 12484 29116 12540
rect 29116 12484 29172 12540
rect 29172 12484 29176 12540
rect 29112 12480 29176 12484
rect 29192 12540 29256 12544
rect 29192 12484 29196 12540
rect 29196 12484 29252 12540
rect 29252 12484 29256 12540
rect 29192 12480 29256 12484
rect 29272 12540 29336 12544
rect 29272 12484 29276 12540
rect 29276 12484 29332 12540
rect 29332 12484 29336 12540
rect 29272 12480 29336 12484
rect 29352 12540 29416 12544
rect 29352 12484 29356 12540
rect 29356 12484 29412 12540
rect 29412 12484 29416 12540
rect 29352 12480 29416 12484
rect 12216 11996 12280 12000
rect 12216 11940 12220 11996
rect 12220 11940 12276 11996
rect 12276 11940 12280 11996
rect 12216 11936 12280 11940
rect 12296 11996 12360 12000
rect 12296 11940 12300 11996
rect 12300 11940 12356 11996
rect 12356 11940 12360 11996
rect 12296 11936 12360 11940
rect 12376 11996 12440 12000
rect 12376 11940 12380 11996
rect 12380 11940 12436 11996
rect 12436 11940 12440 11996
rect 12376 11936 12440 11940
rect 12456 11996 12520 12000
rect 12456 11940 12460 11996
rect 12460 11940 12516 11996
rect 12516 11940 12520 11996
rect 12456 11936 12520 11940
rect 23480 11996 23544 12000
rect 23480 11940 23484 11996
rect 23484 11940 23540 11996
rect 23540 11940 23544 11996
rect 23480 11936 23544 11940
rect 23560 11996 23624 12000
rect 23560 11940 23564 11996
rect 23564 11940 23620 11996
rect 23620 11940 23624 11996
rect 23560 11936 23624 11940
rect 23640 11996 23704 12000
rect 23640 11940 23644 11996
rect 23644 11940 23700 11996
rect 23700 11940 23704 11996
rect 23640 11936 23704 11940
rect 23720 11996 23784 12000
rect 23720 11940 23724 11996
rect 23724 11940 23780 11996
rect 23780 11940 23784 11996
rect 23720 11936 23784 11940
rect 6584 11452 6648 11456
rect 6584 11396 6588 11452
rect 6588 11396 6644 11452
rect 6644 11396 6648 11452
rect 6584 11392 6648 11396
rect 6664 11452 6728 11456
rect 6664 11396 6668 11452
rect 6668 11396 6724 11452
rect 6724 11396 6728 11452
rect 6664 11392 6728 11396
rect 6744 11452 6808 11456
rect 6744 11396 6748 11452
rect 6748 11396 6804 11452
rect 6804 11396 6808 11452
rect 6744 11392 6808 11396
rect 6824 11452 6888 11456
rect 6824 11396 6828 11452
rect 6828 11396 6884 11452
rect 6884 11396 6888 11452
rect 6824 11392 6888 11396
rect 17848 11452 17912 11456
rect 17848 11396 17852 11452
rect 17852 11396 17908 11452
rect 17908 11396 17912 11452
rect 17848 11392 17912 11396
rect 17928 11452 17992 11456
rect 17928 11396 17932 11452
rect 17932 11396 17988 11452
rect 17988 11396 17992 11452
rect 17928 11392 17992 11396
rect 18008 11452 18072 11456
rect 18008 11396 18012 11452
rect 18012 11396 18068 11452
rect 18068 11396 18072 11452
rect 18008 11392 18072 11396
rect 18088 11452 18152 11456
rect 18088 11396 18092 11452
rect 18092 11396 18148 11452
rect 18148 11396 18152 11452
rect 18088 11392 18152 11396
rect 29112 11452 29176 11456
rect 29112 11396 29116 11452
rect 29116 11396 29172 11452
rect 29172 11396 29176 11452
rect 29112 11392 29176 11396
rect 29192 11452 29256 11456
rect 29192 11396 29196 11452
rect 29196 11396 29252 11452
rect 29252 11396 29256 11452
rect 29192 11392 29256 11396
rect 29272 11452 29336 11456
rect 29272 11396 29276 11452
rect 29276 11396 29332 11452
rect 29332 11396 29336 11452
rect 29272 11392 29336 11396
rect 29352 11452 29416 11456
rect 29352 11396 29356 11452
rect 29356 11396 29412 11452
rect 29412 11396 29416 11452
rect 29352 11392 29416 11396
rect 12216 10908 12280 10912
rect 12216 10852 12220 10908
rect 12220 10852 12276 10908
rect 12276 10852 12280 10908
rect 12216 10848 12280 10852
rect 12296 10908 12360 10912
rect 12296 10852 12300 10908
rect 12300 10852 12356 10908
rect 12356 10852 12360 10908
rect 12296 10848 12360 10852
rect 12376 10908 12440 10912
rect 12376 10852 12380 10908
rect 12380 10852 12436 10908
rect 12436 10852 12440 10908
rect 12376 10848 12440 10852
rect 12456 10908 12520 10912
rect 12456 10852 12460 10908
rect 12460 10852 12516 10908
rect 12516 10852 12520 10908
rect 12456 10848 12520 10852
rect 23480 10908 23544 10912
rect 23480 10852 23484 10908
rect 23484 10852 23540 10908
rect 23540 10852 23544 10908
rect 23480 10848 23544 10852
rect 23560 10908 23624 10912
rect 23560 10852 23564 10908
rect 23564 10852 23620 10908
rect 23620 10852 23624 10908
rect 23560 10848 23624 10852
rect 23640 10908 23704 10912
rect 23640 10852 23644 10908
rect 23644 10852 23700 10908
rect 23700 10852 23704 10908
rect 23640 10848 23704 10852
rect 23720 10908 23784 10912
rect 23720 10852 23724 10908
rect 23724 10852 23780 10908
rect 23780 10852 23784 10908
rect 23720 10848 23784 10852
rect 6584 10364 6648 10368
rect 6584 10308 6588 10364
rect 6588 10308 6644 10364
rect 6644 10308 6648 10364
rect 6584 10304 6648 10308
rect 6664 10364 6728 10368
rect 6664 10308 6668 10364
rect 6668 10308 6724 10364
rect 6724 10308 6728 10364
rect 6664 10304 6728 10308
rect 6744 10364 6808 10368
rect 6744 10308 6748 10364
rect 6748 10308 6804 10364
rect 6804 10308 6808 10364
rect 6744 10304 6808 10308
rect 6824 10364 6888 10368
rect 6824 10308 6828 10364
rect 6828 10308 6884 10364
rect 6884 10308 6888 10364
rect 6824 10304 6888 10308
rect 17848 10364 17912 10368
rect 17848 10308 17852 10364
rect 17852 10308 17908 10364
rect 17908 10308 17912 10364
rect 17848 10304 17912 10308
rect 17928 10364 17992 10368
rect 17928 10308 17932 10364
rect 17932 10308 17988 10364
rect 17988 10308 17992 10364
rect 17928 10304 17992 10308
rect 18008 10364 18072 10368
rect 18008 10308 18012 10364
rect 18012 10308 18068 10364
rect 18068 10308 18072 10364
rect 18008 10304 18072 10308
rect 18088 10364 18152 10368
rect 18088 10308 18092 10364
rect 18092 10308 18148 10364
rect 18148 10308 18152 10364
rect 18088 10304 18152 10308
rect 29112 10364 29176 10368
rect 29112 10308 29116 10364
rect 29116 10308 29172 10364
rect 29172 10308 29176 10364
rect 29112 10304 29176 10308
rect 29192 10364 29256 10368
rect 29192 10308 29196 10364
rect 29196 10308 29252 10364
rect 29252 10308 29256 10364
rect 29192 10304 29256 10308
rect 29272 10364 29336 10368
rect 29272 10308 29276 10364
rect 29276 10308 29332 10364
rect 29332 10308 29336 10364
rect 29272 10304 29336 10308
rect 29352 10364 29416 10368
rect 29352 10308 29356 10364
rect 29356 10308 29412 10364
rect 29412 10308 29416 10364
rect 29352 10304 29416 10308
rect 12216 9820 12280 9824
rect 12216 9764 12220 9820
rect 12220 9764 12276 9820
rect 12276 9764 12280 9820
rect 12216 9760 12280 9764
rect 12296 9820 12360 9824
rect 12296 9764 12300 9820
rect 12300 9764 12356 9820
rect 12356 9764 12360 9820
rect 12296 9760 12360 9764
rect 12376 9820 12440 9824
rect 12376 9764 12380 9820
rect 12380 9764 12436 9820
rect 12436 9764 12440 9820
rect 12376 9760 12440 9764
rect 12456 9820 12520 9824
rect 12456 9764 12460 9820
rect 12460 9764 12516 9820
rect 12516 9764 12520 9820
rect 12456 9760 12520 9764
rect 23480 9820 23544 9824
rect 23480 9764 23484 9820
rect 23484 9764 23540 9820
rect 23540 9764 23544 9820
rect 23480 9760 23544 9764
rect 23560 9820 23624 9824
rect 23560 9764 23564 9820
rect 23564 9764 23620 9820
rect 23620 9764 23624 9820
rect 23560 9760 23624 9764
rect 23640 9820 23704 9824
rect 23640 9764 23644 9820
rect 23644 9764 23700 9820
rect 23700 9764 23704 9820
rect 23640 9760 23704 9764
rect 23720 9820 23784 9824
rect 23720 9764 23724 9820
rect 23724 9764 23780 9820
rect 23780 9764 23784 9820
rect 23720 9760 23784 9764
rect 6584 9276 6648 9280
rect 6584 9220 6588 9276
rect 6588 9220 6644 9276
rect 6644 9220 6648 9276
rect 6584 9216 6648 9220
rect 6664 9276 6728 9280
rect 6664 9220 6668 9276
rect 6668 9220 6724 9276
rect 6724 9220 6728 9276
rect 6664 9216 6728 9220
rect 6744 9276 6808 9280
rect 6744 9220 6748 9276
rect 6748 9220 6804 9276
rect 6804 9220 6808 9276
rect 6744 9216 6808 9220
rect 6824 9276 6888 9280
rect 6824 9220 6828 9276
rect 6828 9220 6884 9276
rect 6884 9220 6888 9276
rect 6824 9216 6888 9220
rect 17848 9276 17912 9280
rect 17848 9220 17852 9276
rect 17852 9220 17908 9276
rect 17908 9220 17912 9276
rect 17848 9216 17912 9220
rect 17928 9276 17992 9280
rect 17928 9220 17932 9276
rect 17932 9220 17988 9276
rect 17988 9220 17992 9276
rect 17928 9216 17992 9220
rect 18008 9276 18072 9280
rect 18008 9220 18012 9276
rect 18012 9220 18068 9276
rect 18068 9220 18072 9276
rect 18008 9216 18072 9220
rect 18088 9276 18152 9280
rect 18088 9220 18092 9276
rect 18092 9220 18148 9276
rect 18148 9220 18152 9276
rect 18088 9216 18152 9220
rect 29112 9276 29176 9280
rect 29112 9220 29116 9276
rect 29116 9220 29172 9276
rect 29172 9220 29176 9276
rect 29112 9216 29176 9220
rect 29192 9276 29256 9280
rect 29192 9220 29196 9276
rect 29196 9220 29252 9276
rect 29252 9220 29256 9276
rect 29192 9216 29256 9220
rect 29272 9276 29336 9280
rect 29272 9220 29276 9276
rect 29276 9220 29332 9276
rect 29332 9220 29336 9276
rect 29272 9216 29336 9220
rect 29352 9276 29416 9280
rect 29352 9220 29356 9276
rect 29356 9220 29412 9276
rect 29412 9220 29416 9276
rect 29352 9216 29416 9220
rect 12216 8732 12280 8736
rect 12216 8676 12220 8732
rect 12220 8676 12276 8732
rect 12276 8676 12280 8732
rect 12216 8672 12280 8676
rect 12296 8732 12360 8736
rect 12296 8676 12300 8732
rect 12300 8676 12356 8732
rect 12356 8676 12360 8732
rect 12296 8672 12360 8676
rect 12376 8732 12440 8736
rect 12376 8676 12380 8732
rect 12380 8676 12436 8732
rect 12436 8676 12440 8732
rect 12376 8672 12440 8676
rect 12456 8732 12520 8736
rect 12456 8676 12460 8732
rect 12460 8676 12516 8732
rect 12516 8676 12520 8732
rect 12456 8672 12520 8676
rect 23480 8732 23544 8736
rect 23480 8676 23484 8732
rect 23484 8676 23540 8732
rect 23540 8676 23544 8732
rect 23480 8672 23544 8676
rect 23560 8732 23624 8736
rect 23560 8676 23564 8732
rect 23564 8676 23620 8732
rect 23620 8676 23624 8732
rect 23560 8672 23624 8676
rect 23640 8732 23704 8736
rect 23640 8676 23644 8732
rect 23644 8676 23700 8732
rect 23700 8676 23704 8732
rect 23640 8672 23704 8676
rect 23720 8732 23784 8736
rect 23720 8676 23724 8732
rect 23724 8676 23780 8732
rect 23780 8676 23784 8732
rect 23720 8672 23784 8676
rect 6584 8188 6648 8192
rect 6584 8132 6588 8188
rect 6588 8132 6644 8188
rect 6644 8132 6648 8188
rect 6584 8128 6648 8132
rect 6664 8188 6728 8192
rect 6664 8132 6668 8188
rect 6668 8132 6724 8188
rect 6724 8132 6728 8188
rect 6664 8128 6728 8132
rect 6744 8188 6808 8192
rect 6744 8132 6748 8188
rect 6748 8132 6804 8188
rect 6804 8132 6808 8188
rect 6744 8128 6808 8132
rect 6824 8188 6888 8192
rect 6824 8132 6828 8188
rect 6828 8132 6884 8188
rect 6884 8132 6888 8188
rect 6824 8128 6888 8132
rect 17848 8188 17912 8192
rect 17848 8132 17852 8188
rect 17852 8132 17908 8188
rect 17908 8132 17912 8188
rect 17848 8128 17912 8132
rect 17928 8188 17992 8192
rect 17928 8132 17932 8188
rect 17932 8132 17988 8188
rect 17988 8132 17992 8188
rect 17928 8128 17992 8132
rect 18008 8188 18072 8192
rect 18008 8132 18012 8188
rect 18012 8132 18068 8188
rect 18068 8132 18072 8188
rect 18008 8128 18072 8132
rect 18088 8188 18152 8192
rect 18088 8132 18092 8188
rect 18092 8132 18148 8188
rect 18148 8132 18152 8188
rect 18088 8128 18152 8132
rect 29112 8188 29176 8192
rect 29112 8132 29116 8188
rect 29116 8132 29172 8188
rect 29172 8132 29176 8188
rect 29112 8128 29176 8132
rect 29192 8188 29256 8192
rect 29192 8132 29196 8188
rect 29196 8132 29252 8188
rect 29252 8132 29256 8188
rect 29192 8128 29256 8132
rect 29272 8188 29336 8192
rect 29272 8132 29276 8188
rect 29276 8132 29332 8188
rect 29332 8132 29336 8188
rect 29272 8128 29336 8132
rect 29352 8188 29416 8192
rect 29352 8132 29356 8188
rect 29356 8132 29412 8188
rect 29412 8132 29416 8188
rect 29352 8128 29416 8132
rect 12216 7644 12280 7648
rect 12216 7588 12220 7644
rect 12220 7588 12276 7644
rect 12276 7588 12280 7644
rect 12216 7584 12280 7588
rect 12296 7644 12360 7648
rect 12296 7588 12300 7644
rect 12300 7588 12356 7644
rect 12356 7588 12360 7644
rect 12296 7584 12360 7588
rect 12376 7644 12440 7648
rect 12376 7588 12380 7644
rect 12380 7588 12436 7644
rect 12436 7588 12440 7644
rect 12376 7584 12440 7588
rect 12456 7644 12520 7648
rect 12456 7588 12460 7644
rect 12460 7588 12516 7644
rect 12516 7588 12520 7644
rect 12456 7584 12520 7588
rect 23480 7644 23544 7648
rect 23480 7588 23484 7644
rect 23484 7588 23540 7644
rect 23540 7588 23544 7644
rect 23480 7584 23544 7588
rect 23560 7644 23624 7648
rect 23560 7588 23564 7644
rect 23564 7588 23620 7644
rect 23620 7588 23624 7644
rect 23560 7584 23624 7588
rect 23640 7644 23704 7648
rect 23640 7588 23644 7644
rect 23644 7588 23700 7644
rect 23700 7588 23704 7644
rect 23640 7584 23704 7588
rect 23720 7644 23784 7648
rect 23720 7588 23724 7644
rect 23724 7588 23780 7644
rect 23780 7588 23784 7644
rect 23720 7584 23784 7588
rect 6584 7100 6648 7104
rect 6584 7044 6588 7100
rect 6588 7044 6644 7100
rect 6644 7044 6648 7100
rect 6584 7040 6648 7044
rect 6664 7100 6728 7104
rect 6664 7044 6668 7100
rect 6668 7044 6724 7100
rect 6724 7044 6728 7100
rect 6664 7040 6728 7044
rect 6744 7100 6808 7104
rect 6744 7044 6748 7100
rect 6748 7044 6804 7100
rect 6804 7044 6808 7100
rect 6744 7040 6808 7044
rect 6824 7100 6888 7104
rect 6824 7044 6828 7100
rect 6828 7044 6884 7100
rect 6884 7044 6888 7100
rect 6824 7040 6888 7044
rect 17848 7100 17912 7104
rect 17848 7044 17852 7100
rect 17852 7044 17908 7100
rect 17908 7044 17912 7100
rect 17848 7040 17912 7044
rect 17928 7100 17992 7104
rect 17928 7044 17932 7100
rect 17932 7044 17988 7100
rect 17988 7044 17992 7100
rect 17928 7040 17992 7044
rect 18008 7100 18072 7104
rect 18008 7044 18012 7100
rect 18012 7044 18068 7100
rect 18068 7044 18072 7100
rect 18008 7040 18072 7044
rect 18088 7100 18152 7104
rect 18088 7044 18092 7100
rect 18092 7044 18148 7100
rect 18148 7044 18152 7100
rect 18088 7040 18152 7044
rect 29112 7100 29176 7104
rect 29112 7044 29116 7100
rect 29116 7044 29172 7100
rect 29172 7044 29176 7100
rect 29112 7040 29176 7044
rect 29192 7100 29256 7104
rect 29192 7044 29196 7100
rect 29196 7044 29252 7100
rect 29252 7044 29256 7100
rect 29192 7040 29256 7044
rect 29272 7100 29336 7104
rect 29272 7044 29276 7100
rect 29276 7044 29332 7100
rect 29332 7044 29336 7100
rect 29272 7040 29336 7044
rect 29352 7100 29416 7104
rect 29352 7044 29356 7100
rect 29356 7044 29412 7100
rect 29412 7044 29416 7100
rect 29352 7040 29416 7044
rect 12216 6556 12280 6560
rect 12216 6500 12220 6556
rect 12220 6500 12276 6556
rect 12276 6500 12280 6556
rect 12216 6496 12280 6500
rect 12296 6556 12360 6560
rect 12296 6500 12300 6556
rect 12300 6500 12356 6556
rect 12356 6500 12360 6556
rect 12296 6496 12360 6500
rect 12376 6556 12440 6560
rect 12376 6500 12380 6556
rect 12380 6500 12436 6556
rect 12436 6500 12440 6556
rect 12376 6496 12440 6500
rect 12456 6556 12520 6560
rect 12456 6500 12460 6556
rect 12460 6500 12516 6556
rect 12516 6500 12520 6556
rect 12456 6496 12520 6500
rect 23480 6556 23544 6560
rect 23480 6500 23484 6556
rect 23484 6500 23540 6556
rect 23540 6500 23544 6556
rect 23480 6496 23544 6500
rect 23560 6556 23624 6560
rect 23560 6500 23564 6556
rect 23564 6500 23620 6556
rect 23620 6500 23624 6556
rect 23560 6496 23624 6500
rect 23640 6556 23704 6560
rect 23640 6500 23644 6556
rect 23644 6500 23700 6556
rect 23700 6500 23704 6556
rect 23640 6496 23704 6500
rect 23720 6556 23784 6560
rect 23720 6500 23724 6556
rect 23724 6500 23780 6556
rect 23780 6500 23784 6556
rect 23720 6496 23784 6500
rect 6584 6012 6648 6016
rect 6584 5956 6588 6012
rect 6588 5956 6644 6012
rect 6644 5956 6648 6012
rect 6584 5952 6648 5956
rect 6664 6012 6728 6016
rect 6664 5956 6668 6012
rect 6668 5956 6724 6012
rect 6724 5956 6728 6012
rect 6664 5952 6728 5956
rect 6744 6012 6808 6016
rect 6744 5956 6748 6012
rect 6748 5956 6804 6012
rect 6804 5956 6808 6012
rect 6744 5952 6808 5956
rect 6824 6012 6888 6016
rect 6824 5956 6828 6012
rect 6828 5956 6884 6012
rect 6884 5956 6888 6012
rect 6824 5952 6888 5956
rect 17848 6012 17912 6016
rect 17848 5956 17852 6012
rect 17852 5956 17908 6012
rect 17908 5956 17912 6012
rect 17848 5952 17912 5956
rect 17928 6012 17992 6016
rect 17928 5956 17932 6012
rect 17932 5956 17988 6012
rect 17988 5956 17992 6012
rect 17928 5952 17992 5956
rect 18008 6012 18072 6016
rect 18008 5956 18012 6012
rect 18012 5956 18068 6012
rect 18068 5956 18072 6012
rect 18008 5952 18072 5956
rect 18088 6012 18152 6016
rect 18088 5956 18092 6012
rect 18092 5956 18148 6012
rect 18148 5956 18152 6012
rect 18088 5952 18152 5956
rect 29112 6012 29176 6016
rect 29112 5956 29116 6012
rect 29116 5956 29172 6012
rect 29172 5956 29176 6012
rect 29112 5952 29176 5956
rect 29192 6012 29256 6016
rect 29192 5956 29196 6012
rect 29196 5956 29252 6012
rect 29252 5956 29256 6012
rect 29192 5952 29256 5956
rect 29272 6012 29336 6016
rect 29272 5956 29276 6012
rect 29276 5956 29332 6012
rect 29332 5956 29336 6012
rect 29272 5952 29336 5956
rect 29352 6012 29416 6016
rect 29352 5956 29356 6012
rect 29356 5956 29412 6012
rect 29412 5956 29416 6012
rect 29352 5952 29416 5956
rect 12216 5468 12280 5472
rect 12216 5412 12220 5468
rect 12220 5412 12276 5468
rect 12276 5412 12280 5468
rect 12216 5408 12280 5412
rect 12296 5468 12360 5472
rect 12296 5412 12300 5468
rect 12300 5412 12356 5468
rect 12356 5412 12360 5468
rect 12296 5408 12360 5412
rect 12376 5468 12440 5472
rect 12376 5412 12380 5468
rect 12380 5412 12436 5468
rect 12436 5412 12440 5468
rect 12376 5408 12440 5412
rect 12456 5468 12520 5472
rect 12456 5412 12460 5468
rect 12460 5412 12516 5468
rect 12516 5412 12520 5468
rect 12456 5408 12520 5412
rect 23480 5468 23544 5472
rect 23480 5412 23484 5468
rect 23484 5412 23540 5468
rect 23540 5412 23544 5468
rect 23480 5408 23544 5412
rect 23560 5468 23624 5472
rect 23560 5412 23564 5468
rect 23564 5412 23620 5468
rect 23620 5412 23624 5468
rect 23560 5408 23624 5412
rect 23640 5468 23704 5472
rect 23640 5412 23644 5468
rect 23644 5412 23700 5468
rect 23700 5412 23704 5468
rect 23640 5408 23704 5412
rect 23720 5468 23784 5472
rect 23720 5412 23724 5468
rect 23724 5412 23780 5468
rect 23780 5412 23784 5468
rect 23720 5408 23784 5412
rect 6584 4924 6648 4928
rect 6584 4868 6588 4924
rect 6588 4868 6644 4924
rect 6644 4868 6648 4924
rect 6584 4864 6648 4868
rect 6664 4924 6728 4928
rect 6664 4868 6668 4924
rect 6668 4868 6724 4924
rect 6724 4868 6728 4924
rect 6664 4864 6728 4868
rect 6744 4924 6808 4928
rect 6744 4868 6748 4924
rect 6748 4868 6804 4924
rect 6804 4868 6808 4924
rect 6744 4864 6808 4868
rect 6824 4924 6888 4928
rect 6824 4868 6828 4924
rect 6828 4868 6884 4924
rect 6884 4868 6888 4924
rect 6824 4864 6888 4868
rect 17848 4924 17912 4928
rect 17848 4868 17852 4924
rect 17852 4868 17908 4924
rect 17908 4868 17912 4924
rect 17848 4864 17912 4868
rect 17928 4924 17992 4928
rect 17928 4868 17932 4924
rect 17932 4868 17988 4924
rect 17988 4868 17992 4924
rect 17928 4864 17992 4868
rect 18008 4924 18072 4928
rect 18008 4868 18012 4924
rect 18012 4868 18068 4924
rect 18068 4868 18072 4924
rect 18008 4864 18072 4868
rect 18088 4924 18152 4928
rect 18088 4868 18092 4924
rect 18092 4868 18148 4924
rect 18148 4868 18152 4924
rect 18088 4864 18152 4868
rect 29112 4924 29176 4928
rect 29112 4868 29116 4924
rect 29116 4868 29172 4924
rect 29172 4868 29176 4924
rect 29112 4864 29176 4868
rect 29192 4924 29256 4928
rect 29192 4868 29196 4924
rect 29196 4868 29252 4924
rect 29252 4868 29256 4924
rect 29192 4864 29256 4868
rect 29272 4924 29336 4928
rect 29272 4868 29276 4924
rect 29276 4868 29332 4924
rect 29332 4868 29336 4924
rect 29272 4864 29336 4868
rect 29352 4924 29416 4928
rect 29352 4868 29356 4924
rect 29356 4868 29412 4924
rect 29412 4868 29416 4924
rect 29352 4864 29416 4868
rect 12216 4380 12280 4384
rect 12216 4324 12220 4380
rect 12220 4324 12276 4380
rect 12276 4324 12280 4380
rect 12216 4320 12280 4324
rect 12296 4380 12360 4384
rect 12296 4324 12300 4380
rect 12300 4324 12356 4380
rect 12356 4324 12360 4380
rect 12296 4320 12360 4324
rect 12376 4380 12440 4384
rect 12376 4324 12380 4380
rect 12380 4324 12436 4380
rect 12436 4324 12440 4380
rect 12376 4320 12440 4324
rect 12456 4380 12520 4384
rect 12456 4324 12460 4380
rect 12460 4324 12516 4380
rect 12516 4324 12520 4380
rect 12456 4320 12520 4324
rect 23480 4380 23544 4384
rect 23480 4324 23484 4380
rect 23484 4324 23540 4380
rect 23540 4324 23544 4380
rect 23480 4320 23544 4324
rect 23560 4380 23624 4384
rect 23560 4324 23564 4380
rect 23564 4324 23620 4380
rect 23620 4324 23624 4380
rect 23560 4320 23624 4324
rect 23640 4380 23704 4384
rect 23640 4324 23644 4380
rect 23644 4324 23700 4380
rect 23700 4324 23704 4380
rect 23640 4320 23704 4324
rect 23720 4380 23784 4384
rect 23720 4324 23724 4380
rect 23724 4324 23780 4380
rect 23780 4324 23784 4380
rect 23720 4320 23784 4324
rect 6584 3836 6648 3840
rect 6584 3780 6588 3836
rect 6588 3780 6644 3836
rect 6644 3780 6648 3836
rect 6584 3776 6648 3780
rect 6664 3836 6728 3840
rect 6664 3780 6668 3836
rect 6668 3780 6724 3836
rect 6724 3780 6728 3836
rect 6664 3776 6728 3780
rect 6744 3836 6808 3840
rect 6744 3780 6748 3836
rect 6748 3780 6804 3836
rect 6804 3780 6808 3836
rect 6744 3776 6808 3780
rect 6824 3836 6888 3840
rect 6824 3780 6828 3836
rect 6828 3780 6884 3836
rect 6884 3780 6888 3836
rect 6824 3776 6888 3780
rect 17848 3836 17912 3840
rect 17848 3780 17852 3836
rect 17852 3780 17908 3836
rect 17908 3780 17912 3836
rect 17848 3776 17912 3780
rect 17928 3836 17992 3840
rect 17928 3780 17932 3836
rect 17932 3780 17988 3836
rect 17988 3780 17992 3836
rect 17928 3776 17992 3780
rect 18008 3836 18072 3840
rect 18008 3780 18012 3836
rect 18012 3780 18068 3836
rect 18068 3780 18072 3836
rect 18008 3776 18072 3780
rect 18088 3836 18152 3840
rect 18088 3780 18092 3836
rect 18092 3780 18148 3836
rect 18148 3780 18152 3836
rect 18088 3776 18152 3780
rect 29112 3836 29176 3840
rect 29112 3780 29116 3836
rect 29116 3780 29172 3836
rect 29172 3780 29176 3836
rect 29112 3776 29176 3780
rect 29192 3836 29256 3840
rect 29192 3780 29196 3836
rect 29196 3780 29252 3836
rect 29252 3780 29256 3836
rect 29192 3776 29256 3780
rect 29272 3836 29336 3840
rect 29272 3780 29276 3836
rect 29276 3780 29332 3836
rect 29332 3780 29336 3836
rect 29272 3776 29336 3780
rect 29352 3836 29416 3840
rect 29352 3780 29356 3836
rect 29356 3780 29412 3836
rect 29412 3780 29416 3836
rect 29352 3776 29416 3780
rect 12216 3292 12280 3296
rect 12216 3236 12220 3292
rect 12220 3236 12276 3292
rect 12276 3236 12280 3292
rect 12216 3232 12280 3236
rect 12296 3292 12360 3296
rect 12296 3236 12300 3292
rect 12300 3236 12356 3292
rect 12356 3236 12360 3292
rect 12296 3232 12360 3236
rect 12376 3292 12440 3296
rect 12376 3236 12380 3292
rect 12380 3236 12436 3292
rect 12436 3236 12440 3292
rect 12376 3232 12440 3236
rect 12456 3292 12520 3296
rect 12456 3236 12460 3292
rect 12460 3236 12516 3292
rect 12516 3236 12520 3292
rect 12456 3232 12520 3236
rect 23480 3292 23544 3296
rect 23480 3236 23484 3292
rect 23484 3236 23540 3292
rect 23540 3236 23544 3292
rect 23480 3232 23544 3236
rect 23560 3292 23624 3296
rect 23560 3236 23564 3292
rect 23564 3236 23620 3292
rect 23620 3236 23624 3292
rect 23560 3232 23624 3236
rect 23640 3292 23704 3296
rect 23640 3236 23644 3292
rect 23644 3236 23700 3292
rect 23700 3236 23704 3292
rect 23640 3232 23704 3236
rect 23720 3292 23784 3296
rect 23720 3236 23724 3292
rect 23724 3236 23780 3292
rect 23780 3236 23784 3292
rect 23720 3232 23784 3236
rect 6584 2748 6648 2752
rect 6584 2692 6588 2748
rect 6588 2692 6644 2748
rect 6644 2692 6648 2748
rect 6584 2688 6648 2692
rect 6664 2748 6728 2752
rect 6664 2692 6668 2748
rect 6668 2692 6724 2748
rect 6724 2692 6728 2748
rect 6664 2688 6728 2692
rect 6744 2748 6808 2752
rect 6744 2692 6748 2748
rect 6748 2692 6804 2748
rect 6804 2692 6808 2748
rect 6744 2688 6808 2692
rect 6824 2748 6888 2752
rect 6824 2692 6828 2748
rect 6828 2692 6884 2748
rect 6884 2692 6888 2748
rect 6824 2688 6888 2692
rect 17848 2748 17912 2752
rect 17848 2692 17852 2748
rect 17852 2692 17908 2748
rect 17908 2692 17912 2748
rect 17848 2688 17912 2692
rect 17928 2748 17992 2752
rect 17928 2692 17932 2748
rect 17932 2692 17988 2748
rect 17988 2692 17992 2748
rect 17928 2688 17992 2692
rect 18008 2748 18072 2752
rect 18008 2692 18012 2748
rect 18012 2692 18068 2748
rect 18068 2692 18072 2748
rect 18008 2688 18072 2692
rect 18088 2748 18152 2752
rect 18088 2692 18092 2748
rect 18092 2692 18148 2748
rect 18148 2692 18152 2748
rect 18088 2688 18152 2692
rect 29112 2748 29176 2752
rect 29112 2692 29116 2748
rect 29116 2692 29172 2748
rect 29172 2692 29176 2748
rect 29112 2688 29176 2692
rect 29192 2748 29256 2752
rect 29192 2692 29196 2748
rect 29196 2692 29252 2748
rect 29252 2692 29256 2748
rect 29192 2688 29256 2692
rect 29272 2748 29336 2752
rect 29272 2692 29276 2748
rect 29276 2692 29332 2748
rect 29332 2692 29336 2748
rect 29272 2688 29336 2692
rect 29352 2748 29416 2752
rect 29352 2692 29356 2748
rect 29356 2692 29412 2748
rect 29412 2692 29416 2748
rect 29352 2688 29416 2692
rect 12216 2204 12280 2208
rect 12216 2148 12220 2204
rect 12220 2148 12276 2204
rect 12276 2148 12280 2204
rect 12216 2144 12280 2148
rect 12296 2204 12360 2208
rect 12296 2148 12300 2204
rect 12300 2148 12356 2204
rect 12356 2148 12360 2204
rect 12296 2144 12360 2148
rect 12376 2204 12440 2208
rect 12376 2148 12380 2204
rect 12380 2148 12436 2204
rect 12436 2148 12440 2204
rect 12376 2144 12440 2148
rect 12456 2204 12520 2208
rect 12456 2148 12460 2204
rect 12460 2148 12516 2204
rect 12516 2148 12520 2204
rect 12456 2144 12520 2148
rect 23480 2204 23544 2208
rect 23480 2148 23484 2204
rect 23484 2148 23540 2204
rect 23540 2148 23544 2204
rect 23480 2144 23544 2148
rect 23560 2204 23624 2208
rect 23560 2148 23564 2204
rect 23564 2148 23620 2204
rect 23620 2148 23624 2204
rect 23560 2144 23624 2148
rect 23640 2204 23704 2208
rect 23640 2148 23644 2204
rect 23644 2148 23700 2204
rect 23700 2148 23704 2204
rect 23640 2144 23704 2148
rect 23720 2204 23784 2208
rect 23720 2148 23724 2204
rect 23724 2148 23780 2204
rect 23780 2148 23784 2204
rect 23720 2144 23784 2148
<< metal4 >>
rect 6576 33216 6896 33776
rect 6576 33152 6584 33216
rect 6648 33152 6664 33216
rect 6728 33152 6744 33216
rect 6808 33152 6824 33216
rect 6888 33152 6896 33216
rect 6576 32128 6896 33152
rect 6576 32064 6584 32128
rect 6648 32064 6664 32128
rect 6728 32064 6744 32128
rect 6808 32064 6824 32128
rect 6888 32064 6896 32128
rect 6576 31040 6896 32064
rect 6576 30976 6584 31040
rect 6648 30976 6664 31040
rect 6728 30976 6744 31040
rect 6808 30976 6824 31040
rect 6888 30976 6896 31040
rect 6576 29952 6896 30976
rect 6576 29888 6584 29952
rect 6648 29888 6664 29952
rect 6728 29888 6744 29952
rect 6808 29888 6824 29952
rect 6888 29888 6896 29952
rect 6576 28864 6896 29888
rect 6576 28800 6584 28864
rect 6648 28800 6664 28864
rect 6728 28800 6744 28864
rect 6808 28800 6824 28864
rect 6888 28800 6896 28864
rect 6576 27776 6896 28800
rect 6576 27712 6584 27776
rect 6648 27712 6664 27776
rect 6728 27712 6744 27776
rect 6808 27712 6824 27776
rect 6888 27712 6896 27776
rect 6576 26688 6896 27712
rect 6576 26624 6584 26688
rect 6648 26624 6664 26688
rect 6728 26624 6744 26688
rect 6808 26624 6824 26688
rect 6888 26624 6896 26688
rect 6576 25600 6896 26624
rect 6576 25536 6584 25600
rect 6648 25536 6664 25600
rect 6728 25536 6744 25600
rect 6808 25536 6824 25600
rect 6888 25536 6896 25600
rect 6576 24512 6896 25536
rect 6576 24448 6584 24512
rect 6648 24448 6664 24512
rect 6728 24448 6744 24512
rect 6808 24448 6824 24512
rect 6888 24448 6896 24512
rect 6576 23424 6896 24448
rect 6576 23360 6584 23424
rect 6648 23360 6664 23424
rect 6728 23360 6744 23424
rect 6808 23360 6824 23424
rect 6888 23360 6896 23424
rect 6576 22336 6896 23360
rect 6576 22272 6584 22336
rect 6648 22272 6664 22336
rect 6728 22272 6744 22336
rect 6808 22272 6824 22336
rect 6888 22272 6896 22336
rect 6576 21248 6896 22272
rect 6576 21184 6584 21248
rect 6648 21184 6664 21248
rect 6728 21184 6744 21248
rect 6808 21184 6824 21248
rect 6888 21184 6896 21248
rect 6576 20160 6896 21184
rect 6576 20096 6584 20160
rect 6648 20096 6664 20160
rect 6728 20096 6744 20160
rect 6808 20096 6824 20160
rect 6888 20096 6896 20160
rect 6576 19072 6896 20096
rect 6576 19008 6584 19072
rect 6648 19008 6664 19072
rect 6728 19008 6744 19072
rect 6808 19008 6824 19072
rect 6888 19008 6896 19072
rect 6576 17984 6896 19008
rect 6576 17920 6584 17984
rect 6648 17920 6664 17984
rect 6728 17920 6744 17984
rect 6808 17920 6824 17984
rect 6888 17920 6896 17984
rect 6576 16896 6896 17920
rect 6576 16832 6584 16896
rect 6648 16832 6664 16896
rect 6728 16832 6744 16896
rect 6808 16832 6824 16896
rect 6888 16832 6896 16896
rect 6576 15808 6896 16832
rect 6576 15744 6584 15808
rect 6648 15744 6664 15808
rect 6728 15744 6744 15808
rect 6808 15744 6824 15808
rect 6888 15744 6896 15808
rect 6576 14720 6896 15744
rect 6576 14656 6584 14720
rect 6648 14656 6664 14720
rect 6728 14656 6744 14720
rect 6808 14656 6824 14720
rect 6888 14656 6896 14720
rect 6576 13632 6896 14656
rect 6576 13568 6584 13632
rect 6648 13568 6664 13632
rect 6728 13568 6744 13632
rect 6808 13568 6824 13632
rect 6888 13568 6896 13632
rect 6576 12544 6896 13568
rect 6576 12480 6584 12544
rect 6648 12480 6664 12544
rect 6728 12480 6744 12544
rect 6808 12480 6824 12544
rect 6888 12480 6896 12544
rect 6576 11456 6896 12480
rect 6576 11392 6584 11456
rect 6648 11392 6664 11456
rect 6728 11392 6744 11456
rect 6808 11392 6824 11456
rect 6888 11392 6896 11456
rect 6576 10368 6896 11392
rect 6576 10304 6584 10368
rect 6648 10304 6664 10368
rect 6728 10304 6744 10368
rect 6808 10304 6824 10368
rect 6888 10304 6896 10368
rect 6576 9280 6896 10304
rect 6576 9216 6584 9280
rect 6648 9216 6664 9280
rect 6728 9216 6744 9280
rect 6808 9216 6824 9280
rect 6888 9216 6896 9280
rect 6576 8192 6896 9216
rect 6576 8128 6584 8192
rect 6648 8128 6664 8192
rect 6728 8128 6744 8192
rect 6808 8128 6824 8192
rect 6888 8128 6896 8192
rect 6576 7104 6896 8128
rect 6576 7040 6584 7104
rect 6648 7040 6664 7104
rect 6728 7040 6744 7104
rect 6808 7040 6824 7104
rect 6888 7040 6896 7104
rect 6576 6016 6896 7040
rect 6576 5952 6584 6016
rect 6648 5952 6664 6016
rect 6728 5952 6744 6016
rect 6808 5952 6824 6016
rect 6888 5952 6896 6016
rect 6576 4928 6896 5952
rect 6576 4864 6584 4928
rect 6648 4864 6664 4928
rect 6728 4864 6744 4928
rect 6808 4864 6824 4928
rect 6888 4864 6896 4928
rect 6576 3840 6896 4864
rect 6576 3776 6584 3840
rect 6648 3776 6664 3840
rect 6728 3776 6744 3840
rect 6808 3776 6824 3840
rect 6888 3776 6896 3840
rect 6576 2752 6896 3776
rect 6576 2688 6584 2752
rect 6648 2688 6664 2752
rect 6728 2688 6744 2752
rect 6808 2688 6824 2752
rect 6888 2688 6896 2752
rect 6576 2128 6896 2688
rect 12208 33760 12528 33776
rect 12208 33696 12216 33760
rect 12280 33696 12296 33760
rect 12360 33696 12376 33760
rect 12440 33696 12456 33760
rect 12520 33696 12528 33760
rect 12208 32672 12528 33696
rect 12208 32608 12216 32672
rect 12280 32608 12296 32672
rect 12360 32608 12376 32672
rect 12440 32608 12456 32672
rect 12520 32608 12528 32672
rect 12208 31584 12528 32608
rect 12208 31520 12216 31584
rect 12280 31520 12296 31584
rect 12360 31520 12376 31584
rect 12440 31520 12456 31584
rect 12520 31520 12528 31584
rect 12208 30496 12528 31520
rect 12208 30432 12216 30496
rect 12280 30432 12296 30496
rect 12360 30432 12376 30496
rect 12440 30432 12456 30496
rect 12520 30432 12528 30496
rect 12208 29408 12528 30432
rect 12208 29344 12216 29408
rect 12280 29344 12296 29408
rect 12360 29344 12376 29408
rect 12440 29344 12456 29408
rect 12520 29344 12528 29408
rect 12208 28320 12528 29344
rect 12208 28256 12216 28320
rect 12280 28256 12296 28320
rect 12360 28256 12376 28320
rect 12440 28256 12456 28320
rect 12520 28256 12528 28320
rect 12208 27232 12528 28256
rect 12208 27168 12216 27232
rect 12280 27168 12296 27232
rect 12360 27168 12376 27232
rect 12440 27168 12456 27232
rect 12520 27168 12528 27232
rect 12208 26144 12528 27168
rect 12208 26080 12216 26144
rect 12280 26080 12296 26144
rect 12360 26080 12376 26144
rect 12440 26080 12456 26144
rect 12520 26080 12528 26144
rect 12208 25056 12528 26080
rect 12208 24992 12216 25056
rect 12280 24992 12296 25056
rect 12360 24992 12376 25056
rect 12440 24992 12456 25056
rect 12520 24992 12528 25056
rect 12208 23968 12528 24992
rect 12208 23904 12216 23968
rect 12280 23904 12296 23968
rect 12360 23904 12376 23968
rect 12440 23904 12456 23968
rect 12520 23904 12528 23968
rect 12208 22880 12528 23904
rect 12208 22816 12216 22880
rect 12280 22816 12296 22880
rect 12360 22816 12376 22880
rect 12440 22816 12456 22880
rect 12520 22816 12528 22880
rect 12208 21792 12528 22816
rect 12208 21728 12216 21792
rect 12280 21728 12296 21792
rect 12360 21728 12376 21792
rect 12440 21728 12456 21792
rect 12520 21728 12528 21792
rect 12208 20704 12528 21728
rect 12208 20640 12216 20704
rect 12280 20640 12296 20704
rect 12360 20640 12376 20704
rect 12440 20640 12456 20704
rect 12520 20640 12528 20704
rect 12208 19616 12528 20640
rect 12208 19552 12216 19616
rect 12280 19552 12296 19616
rect 12360 19552 12376 19616
rect 12440 19552 12456 19616
rect 12520 19552 12528 19616
rect 12208 18528 12528 19552
rect 12208 18464 12216 18528
rect 12280 18464 12296 18528
rect 12360 18464 12376 18528
rect 12440 18464 12456 18528
rect 12520 18464 12528 18528
rect 12208 17440 12528 18464
rect 12208 17376 12216 17440
rect 12280 17376 12296 17440
rect 12360 17376 12376 17440
rect 12440 17376 12456 17440
rect 12520 17376 12528 17440
rect 12208 16352 12528 17376
rect 12208 16288 12216 16352
rect 12280 16288 12296 16352
rect 12360 16288 12376 16352
rect 12440 16288 12456 16352
rect 12520 16288 12528 16352
rect 12208 15264 12528 16288
rect 12208 15200 12216 15264
rect 12280 15200 12296 15264
rect 12360 15200 12376 15264
rect 12440 15200 12456 15264
rect 12520 15200 12528 15264
rect 12208 14176 12528 15200
rect 12208 14112 12216 14176
rect 12280 14112 12296 14176
rect 12360 14112 12376 14176
rect 12440 14112 12456 14176
rect 12520 14112 12528 14176
rect 12208 13088 12528 14112
rect 12208 13024 12216 13088
rect 12280 13024 12296 13088
rect 12360 13024 12376 13088
rect 12440 13024 12456 13088
rect 12520 13024 12528 13088
rect 12208 12000 12528 13024
rect 12208 11936 12216 12000
rect 12280 11936 12296 12000
rect 12360 11936 12376 12000
rect 12440 11936 12456 12000
rect 12520 11936 12528 12000
rect 12208 10912 12528 11936
rect 12208 10848 12216 10912
rect 12280 10848 12296 10912
rect 12360 10848 12376 10912
rect 12440 10848 12456 10912
rect 12520 10848 12528 10912
rect 12208 9824 12528 10848
rect 12208 9760 12216 9824
rect 12280 9760 12296 9824
rect 12360 9760 12376 9824
rect 12440 9760 12456 9824
rect 12520 9760 12528 9824
rect 12208 8736 12528 9760
rect 12208 8672 12216 8736
rect 12280 8672 12296 8736
rect 12360 8672 12376 8736
rect 12440 8672 12456 8736
rect 12520 8672 12528 8736
rect 12208 7648 12528 8672
rect 12208 7584 12216 7648
rect 12280 7584 12296 7648
rect 12360 7584 12376 7648
rect 12440 7584 12456 7648
rect 12520 7584 12528 7648
rect 12208 6560 12528 7584
rect 12208 6496 12216 6560
rect 12280 6496 12296 6560
rect 12360 6496 12376 6560
rect 12440 6496 12456 6560
rect 12520 6496 12528 6560
rect 12208 5472 12528 6496
rect 12208 5408 12216 5472
rect 12280 5408 12296 5472
rect 12360 5408 12376 5472
rect 12440 5408 12456 5472
rect 12520 5408 12528 5472
rect 12208 4384 12528 5408
rect 12208 4320 12216 4384
rect 12280 4320 12296 4384
rect 12360 4320 12376 4384
rect 12440 4320 12456 4384
rect 12520 4320 12528 4384
rect 12208 3296 12528 4320
rect 12208 3232 12216 3296
rect 12280 3232 12296 3296
rect 12360 3232 12376 3296
rect 12440 3232 12456 3296
rect 12520 3232 12528 3296
rect 12208 2208 12528 3232
rect 12208 2144 12216 2208
rect 12280 2144 12296 2208
rect 12360 2144 12376 2208
rect 12440 2144 12456 2208
rect 12520 2144 12528 2208
rect 12208 2128 12528 2144
rect 17840 33216 18160 33776
rect 17840 33152 17848 33216
rect 17912 33152 17928 33216
rect 17992 33152 18008 33216
rect 18072 33152 18088 33216
rect 18152 33152 18160 33216
rect 17840 32128 18160 33152
rect 17840 32064 17848 32128
rect 17912 32064 17928 32128
rect 17992 32064 18008 32128
rect 18072 32064 18088 32128
rect 18152 32064 18160 32128
rect 17840 31040 18160 32064
rect 17840 30976 17848 31040
rect 17912 30976 17928 31040
rect 17992 30976 18008 31040
rect 18072 30976 18088 31040
rect 18152 30976 18160 31040
rect 17840 29952 18160 30976
rect 17840 29888 17848 29952
rect 17912 29888 17928 29952
rect 17992 29888 18008 29952
rect 18072 29888 18088 29952
rect 18152 29888 18160 29952
rect 17840 28864 18160 29888
rect 17840 28800 17848 28864
rect 17912 28800 17928 28864
rect 17992 28800 18008 28864
rect 18072 28800 18088 28864
rect 18152 28800 18160 28864
rect 17840 27776 18160 28800
rect 17840 27712 17848 27776
rect 17912 27712 17928 27776
rect 17992 27712 18008 27776
rect 18072 27712 18088 27776
rect 18152 27712 18160 27776
rect 17840 26688 18160 27712
rect 17840 26624 17848 26688
rect 17912 26624 17928 26688
rect 17992 26624 18008 26688
rect 18072 26624 18088 26688
rect 18152 26624 18160 26688
rect 17840 25600 18160 26624
rect 17840 25536 17848 25600
rect 17912 25536 17928 25600
rect 17992 25536 18008 25600
rect 18072 25536 18088 25600
rect 18152 25536 18160 25600
rect 17840 24512 18160 25536
rect 17840 24448 17848 24512
rect 17912 24448 17928 24512
rect 17992 24448 18008 24512
rect 18072 24448 18088 24512
rect 18152 24448 18160 24512
rect 17840 23424 18160 24448
rect 17840 23360 17848 23424
rect 17912 23360 17928 23424
rect 17992 23360 18008 23424
rect 18072 23360 18088 23424
rect 18152 23360 18160 23424
rect 17840 22336 18160 23360
rect 17840 22272 17848 22336
rect 17912 22272 17928 22336
rect 17992 22272 18008 22336
rect 18072 22272 18088 22336
rect 18152 22272 18160 22336
rect 17840 21248 18160 22272
rect 17840 21184 17848 21248
rect 17912 21184 17928 21248
rect 17992 21184 18008 21248
rect 18072 21184 18088 21248
rect 18152 21184 18160 21248
rect 17840 20160 18160 21184
rect 17840 20096 17848 20160
rect 17912 20096 17928 20160
rect 17992 20096 18008 20160
rect 18072 20096 18088 20160
rect 18152 20096 18160 20160
rect 17840 19072 18160 20096
rect 17840 19008 17848 19072
rect 17912 19008 17928 19072
rect 17992 19008 18008 19072
rect 18072 19008 18088 19072
rect 18152 19008 18160 19072
rect 17840 17984 18160 19008
rect 17840 17920 17848 17984
rect 17912 17920 17928 17984
rect 17992 17920 18008 17984
rect 18072 17920 18088 17984
rect 18152 17920 18160 17984
rect 17840 16896 18160 17920
rect 17840 16832 17848 16896
rect 17912 16832 17928 16896
rect 17992 16832 18008 16896
rect 18072 16832 18088 16896
rect 18152 16832 18160 16896
rect 17840 15808 18160 16832
rect 17840 15744 17848 15808
rect 17912 15744 17928 15808
rect 17992 15744 18008 15808
rect 18072 15744 18088 15808
rect 18152 15744 18160 15808
rect 17840 14720 18160 15744
rect 17840 14656 17848 14720
rect 17912 14656 17928 14720
rect 17992 14656 18008 14720
rect 18072 14656 18088 14720
rect 18152 14656 18160 14720
rect 17840 13632 18160 14656
rect 17840 13568 17848 13632
rect 17912 13568 17928 13632
rect 17992 13568 18008 13632
rect 18072 13568 18088 13632
rect 18152 13568 18160 13632
rect 17840 12544 18160 13568
rect 17840 12480 17848 12544
rect 17912 12480 17928 12544
rect 17992 12480 18008 12544
rect 18072 12480 18088 12544
rect 18152 12480 18160 12544
rect 17840 11456 18160 12480
rect 17840 11392 17848 11456
rect 17912 11392 17928 11456
rect 17992 11392 18008 11456
rect 18072 11392 18088 11456
rect 18152 11392 18160 11456
rect 17840 10368 18160 11392
rect 17840 10304 17848 10368
rect 17912 10304 17928 10368
rect 17992 10304 18008 10368
rect 18072 10304 18088 10368
rect 18152 10304 18160 10368
rect 17840 9280 18160 10304
rect 17840 9216 17848 9280
rect 17912 9216 17928 9280
rect 17992 9216 18008 9280
rect 18072 9216 18088 9280
rect 18152 9216 18160 9280
rect 17840 8192 18160 9216
rect 17840 8128 17848 8192
rect 17912 8128 17928 8192
rect 17992 8128 18008 8192
rect 18072 8128 18088 8192
rect 18152 8128 18160 8192
rect 17840 7104 18160 8128
rect 17840 7040 17848 7104
rect 17912 7040 17928 7104
rect 17992 7040 18008 7104
rect 18072 7040 18088 7104
rect 18152 7040 18160 7104
rect 17840 6016 18160 7040
rect 17840 5952 17848 6016
rect 17912 5952 17928 6016
rect 17992 5952 18008 6016
rect 18072 5952 18088 6016
rect 18152 5952 18160 6016
rect 17840 4928 18160 5952
rect 17840 4864 17848 4928
rect 17912 4864 17928 4928
rect 17992 4864 18008 4928
rect 18072 4864 18088 4928
rect 18152 4864 18160 4928
rect 17840 3840 18160 4864
rect 17840 3776 17848 3840
rect 17912 3776 17928 3840
rect 17992 3776 18008 3840
rect 18072 3776 18088 3840
rect 18152 3776 18160 3840
rect 17840 2752 18160 3776
rect 17840 2688 17848 2752
rect 17912 2688 17928 2752
rect 17992 2688 18008 2752
rect 18072 2688 18088 2752
rect 18152 2688 18160 2752
rect 17840 2128 18160 2688
rect 23472 33760 23792 33776
rect 23472 33696 23480 33760
rect 23544 33696 23560 33760
rect 23624 33696 23640 33760
rect 23704 33696 23720 33760
rect 23784 33696 23792 33760
rect 23472 32672 23792 33696
rect 23472 32608 23480 32672
rect 23544 32608 23560 32672
rect 23624 32608 23640 32672
rect 23704 32608 23720 32672
rect 23784 32608 23792 32672
rect 23472 31584 23792 32608
rect 23472 31520 23480 31584
rect 23544 31520 23560 31584
rect 23624 31520 23640 31584
rect 23704 31520 23720 31584
rect 23784 31520 23792 31584
rect 23472 30496 23792 31520
rect 23472 30432 23480 30496
rect 23544 30432 23560 30496
rect 23624 30432 23640 30496
rect 23704 30432 23720 30496
rect 23784 30432 23792 30496
rect 23472 29408 23792 30432
rect 23472 29344 23480 29408
rect 23544 29344 23560 29408
rect 23624 29344 23640 29408
rect 23704 29344 23720 29408
rect 23784 29344 23792 29408
rect 23472 28320 23792 29344
rect 23472 28256 23480 28320
rect 23544 28256 23560 28320
rect 23624 28256 23640 28320
rect 23704 28256 23720 28320
rect 23784 28256 23792 28320
rect 23472 27232 23792 28256
rect 23472 27168 23480 27232
rect 23544 27168 23560 27232
rect 23624 27168 23640 27232
rect 23704 27168 23720 27232
rect 23784 27168 23792 27232
rect 23472 26144 23792 27168
rect 23472 26080 23480 26144
rect 23544 26080 23560 26144
rect 23624 26080 23640 26144
rect 23704 26080 23720 26144
rect 23784 26080 23792 26144
rect 23472 25056 23792 26080
rect 23472 24992 23480 25056
rect 23544 24992 23560 25056
rect 23624 24992 23640 25056
rect 23704 24992 23720 25056
rect 23784 24992 23792 25056
rect 23472 23968 23792 24992
rect 23472 23904 23480 23968
rect 23544 23904 23560 23968
rect 23624 23904 23640 23968
rect 23704 23904 23720 23968
rect 23784 23904 23792 23968
rect 23472 22880 23792 23904
rect 23472 22816 23480 22880
rect 23544 22816 23560 22880
rect 23624 22816 23640 22880
rect 23704 22816 23720 22880
rect 23784 22816 23792 22880
rect 23472 21792 23792 22816
rect 23472 21728 23480 21792
rect 23544 21728 23560 21792
rect 23624 21728 23640 21792
rect 23704 21728 23720 21792
rect 23784 21728 23792 21792
rect 23472 20704 23792 21728
rect 23472 20640 23480 20704
rect 23544 20640 23560 20704
rect 23624 20640 23640 20704
rect 23704 20640 23720 20704
rect 23784 20640 23792 20704
rect 23472 19616 23792 20640
rect 23472 19552 23480 19616
rect 23544 19552 23560 19616
rect 23624 19552 23640 19616
rect 23704 19552 23720 19616
rect 23784 19552 23792 19616
rect 23472 18528 23792 19552
rect 23472 18464 23480 18528
rect 23544 18464 23560 18528
rect 23624 18464 23640 18528
rect 23704 18464 23720 18528
rect 23784 18464 23792 18528
rect 23472 17440 23792 18464
rect 23472 17376 23480 17440
rect 23544 17376 23560 17440
rect 23624 17376 23640 17440
rect 23704 17376 23720 17440
rect 23784 17376 23792 17440
rect 23472 16352 23792 17376
rect 23472 16288 23480 16352
rect 23544 16288 23560 16352
rect 23624 16288 23640 16352
rect 23704 16288 23720 16352
rect 23784 16288 23792 16352
rect 23472 15264 23792 16288
rect 23472 15200 23480 15264
rect 23544 15200 23560 15264
rect 23624 15200 23640 15264
rect 23704 15200 23720 15264
rect 23784 15200 23792 15264
rect 23472 14176 23792 15200
rect 23472 14112 23480 14176
rect 23544 14112 23560 14176
rect 23624 14112 23640 14176
rect 23704 14112 23720 14176
rect 23784 14112 23792 14176
rect 23472 13088 23792 14112
rect 23472 13024 23480 13088
rect 23544 13024 23560 13088
rect 23624 13024 23640 13088
rect 23704 13024 23720 13088
rect 23784 13024 23792 13088
rect 23472 12000 23792 13024
rect 23472 11936 23480 12000
rect 23544 11936 23560 12000
rect 23624 11936 23640 12000
rect 23704 11936 23720 12000
rect 23784 11936 23792 12000
rect 23472 10912 23792 11936
rect 23472 10848 23480 10912
rect 23544 10848 23560 10912
rect 23624 10848 23640 10912
rect 23704 10848 23720 10912
rect 23784 10848 23792 10912
rect 23472 9824 23792 10848
rect 23472 9760 23480 9824
rect 23544 9760 23560 9824
rect 23624 9760 23640 9824
rect 23704 9760 23720 9824
rect 23784 9760 23792 9824
rect 23472 8736 23792 9760
rect 23472 8672 23480 8736
rect 23544 8672 23560 8736
rect 23624 8672 23640 8736
rect 23704 8672 23720 8736
rect 23784 8672 23792 8736
rect 23472 7648 23792 8672
rect 23472 7584 23480 7648
rect 23544 7584 23560 7648
rect 23624 7584 23640 7648
rect 23704 7584 23720 7648
rect 23784 7584 23792 7648
rect 23472 6560 23792 7584
rect 23472 6496 23480 6560
rect 23544 6496 23560 6560
rect 23624 6496 23640 6560
rect 23704 6496 23720 6560
rect 23784 6496 23792 6560
rect 23472 5472 23792 6496
rect 23472 5408 23480 5472
rect 23544 5408 23560 5472
rect 23624 5408 23640 5472
rect 23704 5408 23720 5472
rect 23784 5408 23792 5472
rect 23472 4384 23792 5408
rect 23472 4320 23480 4384
rect 23544 4320 23560 4384
rect 23624 4320 23640 4384
rect 23704 4320 23720 4384
rect 23784 4320 23792 4384
rect 23472 3296 23792 4320
rect 23472 3232 23480 3296
rect 23544 3232 23560 3296
rect 23624 3232 23640 3296
rect 23704 3232 23720 3296
rect 23784 3232 23792 3296
rect 23472 2208 23792 3232
rect 23472 2144 23480 2208
rect 23544 2144 23560 2208
rect 23624 2144 23640 2208
rect 23704 2144 23720 2208
rect 23784 2144 23792 2208
rect 23472 2128 23792 2144
rect 29104 33216 29424 33776
rect 29104 33152 29112 33216
rect 29176 33152 29192 33216
rect 29256 33152 29272 33216
rect 29336 33152 29352 33216
rect 29416 33152 29424 33216
rect 29104 32128 29424 33152
rect 29104 32064 29112 32128
rect 29176 32064 29192 32128
rect 29256 32064 29272 32128
rect 29336 32064 29352 32128
rect 29416 32064 29424 32128
rect 29104 31040 29424 32064
rect 29104 30976 29112 31040
rect 29176 30976 29192 31040
rect 29256 30976 29272 31040
rect 29336 30976 29352 31040
rect 29416 30976 29424 31040
rect 29104 29952 29424 30976
rect 29104 29888 29112 29952
rect 29176 29888 29192 29952
rect 29256 29888 29272 29952
rect 29336 29888 29352 29952
rect 29416 29888 29424 29952
rect 29104 28864 29424 29888
rect 29104 28800 29112 28864
rect 29176 28800 29192 28864
rect 29256 28800 29272 28864
rect 29336 28800 29352 28864
rect 29416 28800 29424 28864
rect 29104 27776 29424 28800
rect 29104 27712 29112 27776
rect 29176 27712 29192 27776
rect 29256 27712 29272 27776
rect 29336 27712 29352 27776
rect 29416 27712 29424 27776
rect 29104 26688 29424 27712
rect 29104 26624 29112 26688
rect 29176 26624 29192 26688
rect 29256 26624 29272 26688
rect 29336 26624 29352 26688
rect 29416 26624 29424 26688
rect 29104 25600 29424 26624
rect 29104 25536 29112 25600
rect 29176 25536 29192 25600
rect 29256 25536 29272 25600
rect 29336 25536 29352 25600
rect 29416 25536 29424 25600
rect 29104 24512 29424 25536
rect 29104 24448 29112 24512
rect 29176 24448 29192 24512
rect 29256 24448 29272 24512
rect 29336 24448 29352 24512
rect 29416 24448 29424 24512
rect 29104 23424 29424 24448
rect 29104 23360 29112 23424
rect 29176 23360 29192 23424
rect 29256 23360 29272 23424
rect 29336 23360 29352 23424
rect 29416 23360 29424 23424
rect 29104 22336 29424 23360
rect 29104 22272 29112 22336
rect 29176 22272 29192 22336
rect 29256 22272 29272 22336
rect 29336 22272 29352 22336
rect 29416 22272 29424 22336
rect 29104 21248 29424 22272
rect 29104 21184 29112 21248
rect 29176 21184 29192 21248
rect 29256 21184 29272 21248
rect 29336 21184 29352 21248
rect 29416 21184 29424 21248
rect 29104 20160 29424 21184
rect 29104 20096 29112 20160
rect 29176 20096 29192 20160
rect 29256 20096 29272 20160
rect 29336 20096 29352 20160
rect 29416 20096 29424 20160
rect 29104 19072 29424 20096
rect 29104 19008 29112 19072
rect 29176 19008 29192 19072
rect 29256 19008 29272 19072
rect 29336 19008 29352 19072
rect 29416 19008 29424 19072
rect 29104 17984 29424 19008
rect 29104 17920 29112 17984
rect 29176 17920 29192 17984
rect 29256 17920 29272 17984
rect 29336 17920 29352 17984
rect 29416 17920 29424 17984
rect 29104 16896 29424 17920
rect 29104 16832 29112 16896
rect 29176 16832 29192 16896
rect 29256 16832 29272 16896
rect 29336 16832 29352 16896
rect 29416 16832 29424 16896
rect 29104 15808 29424 16832
rect 29104 15744 29112 15808
rect 29176 15744 29192 15808
rect 29256 15744 29272 15808
rect 29336 15744 29352 15808
rect 29416 15744 29424 15808
rect 29104 14720 29424 15744
rect 29104 14656 29112 14720
rect 29176 14656 29192 14720
rect 29256 14656 29272 14720
rect 29336 14656 29352 14720
rect 29416 14656 29424 14720
rect 29104 13632 29424 14656
rect 29104 13568 29112 13632
rect 29176 13568 29192 13632
rect 29256 13568 29272 13632
rect 29336 13568 29352 13632
rect 29416 13568 29424 13632
rect 29104 12544 29424 13568
rect 29104 12480 29112 12544
rect 29176 12480 29192 12544
rect 29256 12480 29272 12544
rect 29336 12480 29352 12544
rect 29416 12480 29424 12544
rect 29104 11456 29424 12480
rect 29104 11392 29112 11456
rect 29176 11392 29192 11456
rect 29256 11392 29272 11456
rect 29336 11392 29352 11456
rect 29416 11392 29424 11456
rect 29104 10368 29424 11392
rect 29104 10304 29112 10368
rect 29176 10304 29192 10368
rect 29256 10304 29272 10368
rect 29336 10304 29352 10368
rect 29416 10304 29424 10368
rect 29104 9280 29424 10304
rect 29104 9216 29112 9280
rect 29176 9216 29192 9280
rect 29256 9216 29272 9280
rect 29336 9216 29352 9280
rect 29416 9216 29424 9280
rect 29104 8192 29424 9216
rect 29104 8128 29112 8192
rect 29176 8128 29192 8192
rect 29256 8128 29272 8192
rect 29336 8128 29352 8192
rect 29416 8128 29424 8192
rect 29104 7104 29424 8128
rect 29104 7040 29112 7104
rect 29176 7040 29192 7104
rect 29256 7040 29272 7104
rect 29336 7040 29352 7104
rect 29416 7040 29424 7104
rect 29104 6016 29424 7040
rect 29104 5952 29112 6016
rect 29176 5952 29192 6016
rect 29256 5952 29272 6016
rect 29336 5952 29352 6016
rect 29416 5952 29424 6016
rect 29104 4928 29424 5952
rect 29104 4864 29112 4928
rect 29176 4864 29192 4928
rect 29256 4864 29272 4928
rect 29336 4864 29352 4928
rect 29416 4864 29424 4928
rect 29104 3840 29424 4864
rect 29104 3776 29112 3840
rect 29176 3776 29192 3840
rect 29256 3776 29272 3840
rect 29336 3776 29352 3840
rect 29416 3776 29424 3840
rect 29104 2752 29424 3776
rect 29104 2688 29112 2752
rect 29176 2688 29192 2752
rect 29256 2688 29272 2752
rect 29336 2688 29352 2752
rect 29416 2688 29424 2752
rect 29104 2128 29424 2688
use sky130_fd_sc_hd__diode_2  ANTENNA__011__A pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 18952 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__012__A
timestamp 1644511149
transform -1 0 21068 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__012__B
timestamp 1644511149
transform -1 0 21988 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__013__B
timestamp 1644511149
transform 1 0 20976 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__014__A
timestamp 1644511149
transform 1 0 20240 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__014__B
timestamp 1644511149
transform 1 0 21252 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__015__B1
timestamp 1644511149
transform 1 0 21896 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__016__C1
timestamp 1644511149
transform 1 0 18860 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__017__A
timestamp 1644511149
transform -1 0 21988 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__019__A
timestamp 1644511149
transform -1 0 21804 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__019__B
timestamp 1644511149
transform 1 0 22172 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__020__A1
timestamp 1644511149
transform 1 0 19228 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__021__A
timestamp 1644511149
transform 1 0 20332 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__022__B1_N
timestamp 1644511149
transform -1 0 19872 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__023__A
timestamp 1644511149
transform -1 0 18676 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__024__B1_N
timestamp 1644511149
transform 1 0 18584 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__027__A
timestamp 1644511149
transform 1 0 16928 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__029__A
timestamp 1644511149
transform -1 0 19412 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__030__A
timestamp 1644511149
transform -1 0 17572 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__032__A
timestamp 1644511149
transform 1 0 16928 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__035__A
timestamp 1644511149
transform -1 0 16376 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__039__A
timestamp 1644511149
transform -1 0 20148 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__040__A
timestamp 1644511149
transform 1 0 18860 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__043__A
timestamp 1644511149
transform 1 0 18400 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__049__A
timestamp 1644511149
transform 1 0 30360 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__050__A
timestamp 1644511149
transform -1 0 16744 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__060__A
timestamp 1644511149
transform 1 0 21160 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__061__A
timestamp 1644511149
transform 1 0 33580 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__076__A
timestamp 1644511149
transform 1 0 18952 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__078__A
timestamp 1644511149
transform -1 0 30452 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__083__A
timestamp 1644511149
transform 1 0 17112 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__084__A
timestamp 1644511149
transform 1 0 17572 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__091__A
timestamp 1644511149
transform -1 0 19136 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__093__A
timestamp 1644511149
transform -1 0 18308 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__105__A
timestamp 1644511149
transform -1 0 19136 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__106__A
timestamp 1644511149
transform 1 0 16008 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1644511149
transform -1 0 2116 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1644511149
transform -1 0 23920 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1644511149
transform -1 0 12328 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1644511149
transform -1 0 34408 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1644511149
transform -1 0 2024 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1644511149
transform -1 0 17572 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1644511149
transform -1 0 3956 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1644511149
transform -1 0 33856 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1644511149
transform -1 0 4876 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1644511149
transform -1 0 33948 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1644511149
transform -1 0 31372 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1644511149
transform -1 0 1564 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1644511149
transform -1 0 33948 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1644511149
transform -1 0 19412 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1644511149
transform -1 0 11684 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1644511149
transform -1 0 30360 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1644511149
transform -1 0 33856 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1644511149
transform -1 0 32844 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1644511149
transform -1 0 3404 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1644511149
transform -1 0 33948 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1644511149
transform -1 0 31832 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1644511149
transform -1 0 5704 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1644511149
transform -1 0 33856 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1644511149
transform -1 0 15916 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1644511149
transform -1 0 2484 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1644511149
transform -1 0 28244 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1644511149
transform -1 0 33948 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1644511149
transform -1 0 12236 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1644511149
transform -1 0 2116 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1644511149
transform -1 0 9752 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1644511149
transform -1 0 30820 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1644511149
transform -1 0 33948 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1644511149
transform -1 0 1564 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1644511149
transform -1 0 24104 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1644511149
transform -1 0 34408 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1644511149
transform -1 0 2024 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1644511149
transform -1 0 2852 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1644511149
transform -1 0 2024 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1644511149
transform -1 0 29256 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1644511149
transform -1 0 2576 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1644511149
transform -1 0 33396 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1644511149
transform -1 0 10856 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1644511149
transform -1 0 3220 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1644511149
transform -1 0 3588 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1644511149
transform -1 0 26680 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1644511149
transform -1 0 33304 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 1644511149
transform -1 0 13432 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 1644511149
transform -1 0 33856 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 1644511149
transform -1 0 30360 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 1644511149
transform -1 0 22632 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input51_A
timestamp 1644511149
transform -1 0 33948 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input52_A
timestamp 1644511149
transform -1 0 2300 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input53_A
timestamp 1644511149
transform -1 0 2300 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input54_A
timestamp 1644511149
transform -1 0 22448 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input55_A
timestamp 1644511149
transform -1 0 29532 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input56_A
timestamp 1644511149
transform -1 0 33028 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input57_A
timestamp 1644511149
transform -1 0 14812 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input58_A
timestamp 1644511149
transform -1 0 1564 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input59_A
timestamp 1644511149
transform -1 0 33948 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input60_A
timestamp 1644511149
transform -1 0 3220 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input61_A
timestamp 1644511149
transform -1 0 33948 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input62_A
timestamp 1644511149
transform -1 0 9292 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input63_A
timestamp 1644511149
transform -1 0 33304 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input64_A
timestamp 1644511149
transform -1 0 32936 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input65_A
timestamp 1644511149
transform -1 0 4600 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input66_A
timestamp 1644511149
transform -1 0 34040 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input67_A
timestamp 1644511149
transform -1 0 19780 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input68_A
timestamp 1644511149
transform -1 0 8464 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input69_A
timestamp 1644511149
transform -1 0 15272 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input70_A
timestamp 1644511149
transform -1 0 26680 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input71_A
timestamp 1644511149
transform -1 0 31832 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input72_A
timestamp 1644511149
transform -1 0 32476 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input73_A
timestamp 1644511149
transform -1 0 33580 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input74_A
timestamp 1644511149
transform -1 0 14720 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input75_A
timestamp 1644511149
transform -1 0 21712 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input76_A
timestamp 1644511149
transform -1 0 18952 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input77_A
timestamp 1644511149
transform -1 0 1564 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input78_A
timestamp 1644511149
transform -1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input79_A
timestamp 1644511149
transform -1 0 33856 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input80_A
timestamp 1644511149
transform -1 0 15548 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input81_A
timestamp 1644511149
transform -1 0 33580 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input82_A
timestamp 1644511149
transform -1 0 8556 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input83_A
timestamp 1644511149
transform -1 0 23092 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input84_A
timestamp 1644511149
transform -1 0 2668 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input85_A
timestamp 1644511149
transform -1 0 33948 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input86_A
timestamp 1644511149
transform -1 0 3128 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input87_A
timestamp 1644511149
transform -1 0 8648 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input88_A
timestamp 1644511149
transform -1 0 34408 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output89_A
timestamp 1644511149
transform 1 0 33396 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output92_A
timestamp 1644511149
transform -1 0 23000 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output95_A
timestamp 1644511149
transform 1 0 1932 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output96_A
timestamp 1644511149
transform 1 0 1932 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output99_A
timestamp 1644511149
transform 1 0 31648 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output107_A
timestamp 1644511149
transform 1 0 4140 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output109_A
timestamp 1644511149
transform 1 0 32384 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output111_A
timestamp 1644511149
transform -1 0 13800 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output114_A
timestamp 1644511149
transform -1 0 27876 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output116_A
timestamp 1644511149
transform 1 0 33672 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output119_A
timestamp 1644511149
transform 1 0 33672 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output122_A
timestamp 1644511149
transform 1 0 31280 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output124_A
timestamp 1644511149
transform -1 0 34040 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output126_A
timestamp 1644511149
transform 1 0 8096 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output127_A
timestamp 1644511149
transform -1 0 33856 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output129_A
timestamp 1644511149
transform -1 0 33488 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output135_A
timestamp 1644511149
transform 1 0 32476 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output136_A
timestamp 1644511149
transform 1 0 33672 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output139_A
timestamp 1644511149
transform -1 0 33856 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output146_A
timestamp 1644511149
transform 1 0 1932 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output150_A
timestamp 1644511149
transform 1 0 1932 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output159_A
timestamp 1644511149
transform 1 0 28704 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output161_A
timestamp 1644511149
transform -1 0 2484 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output165_A
timestamp 1644511149
transform 1 0 1932 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output167_A
timestamp 1644511149
transform -1 0 21068 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output168_A
timestamp 1644511149
transform 1 0 25484 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output170_A
timestamp 1644511149
transform -1 0 3036 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output171_A
timestamp 1644511149
transform -1 0 6624 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output172_A
timestamp 1644511149
transform -1 0 25300 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output173_A
timestamp 1644511149
transform 1 0 1932 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output174_A
timestamp 1644511149
transform -1 0 2116 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2300 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19
timestamp 1644511149
transform 1 0 2852 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3404 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39
timestamp 1644511149
transform 1 0 4692 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 5796 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_67
timestamp 1644511149
transform 1 0 7268 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_73
timestamp 1644511149
transform 1 0 7820 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77
timestamp 1644511149
transform 1 0 8188 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82
timestamp 1644511149
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1644511149
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_97
timestamp 1644511149
transform 1 0 10028 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_103
timestamp 1644511149
transform 1 0 10580 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1644511149
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_113
timestamp 1644511149
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_119
timestamp 1644511149
transform 1 0 12052 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_126
timestamp 1644511149
transform 1 0 12696 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_138
timestamp 1644511149
transform 1 0 13800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_141
timestamp 1644511149
transform 1 0 14076 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_147
timestamp 1644511149
transform 1 0 14628 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_153
timestamp 1644511149
transform 1 0 15180 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_157
timestamp 1644511149
transform 1 0 15548 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_161
timestamp 1644511149
transform 1 0 15916 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_166
timestamp 1644511149
transform 1 0 16376 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_173
timestamp 1644511149
transform 1 0 17020 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_177
timestamp 1644511149
transform 1 0 17388 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_182
timestamp 1644511149
transform 1 0 17848 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_194
timestamp 1644511149
transform 1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_207
timestamp 1644511149
transform 1 0 20148 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_213
timestamp 1644511149
transform 1 0 20700 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_217 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21068 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_223
timestamp 1644511149
transform 1 0 21620 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_229
timestamp 1644511149
transform 1 0 22172 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_233
timestamp 1644511149
transform 1 0 22540 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_238
timestamp 1644511149
transform 1 0 23000 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_244
timestamp 1644511149
transform 1 0 23552 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_248
timestamp 1644511149
transform 1 0 23920 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_257
timestamp 1644511149
transform 1 0 24748 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_261
timestamp 1644511149
transform 1 0 25116 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_266 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25576 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_274
timestamp 1644511149
transform 1 0 26312 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_278
timestamp 1644511149
transform 1 0 26680 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_291
timestamp 1644511149
transform 1 0 27876 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_297
timestamp 1644511149
transform 1 0 28428 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_302
timestamp 1644511149
transform 1 0 28888 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_306
timestamp 1644511149
transform 1 0 29256 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_319
timestamp 1644511149
transform 1 0 30452 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_325
timestamp 1644511149
transform 1 0 31004 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_329
timestamp 1644511149
transform 1 0 31372 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_334
timestamp 1644511149
transform 1 0 31832 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_337
timestamp 1644511149
transform 1 0 32108 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_344
timestamp 1644511149
transform 1 0 32752 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_350
timestamp 1644511149
transform 1 0 33304 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_362
timestamp 1644511149
transform 1 0 34408 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_13
timestamp 1644511149
transform 1 0 2300 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_19
timestamp 1644511149
transform 1 0 2852 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_23
timestamp 1644511149
transform 1 0 3220 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_27
timestamp 1644511149
transform 1 0 3588 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_35
timestamp 1644511149
transform 1 0 4324 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_41
timestamp 1644511149
transform 1 0 4876 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_49
timestamp 1644511149
transform 1 0 5612 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp 1644511149
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_57
timestamp 1644511149
transform 1 0 6348 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_63
timestamp 1644511149
transform 1 0 6900 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_71
timestamp 1644511149
transform 1 0 7636 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_76
timestamp 1644511149
transform 1 0 8096 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_80
timestamp 1644511149
transform 1 0 8464 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_85
timestamp 1644511149
transform 1 0 8924 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_89 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 9292 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_101
timestamp 1644511149
transform 1 0 10396 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_109
timestamp 1644511149
transform 1 0 11132 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_113
timestamp 1644511149
transform 1 0 11500 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_117
timestamp 1644511149
transform 1 0 11868 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_121
timestamp 1644511149
transform 1 0 12236 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_129
timestamp 1644511149
transform 1 0 12972 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_134
timestamp 1644511149
transform 1 0 13432 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_139
timestamp 1644511149
transform 1 0 13892 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_145
timestamp 1644511149
transform 1 0 14444 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_149
timestamp 1644511149
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1644511149
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1644511149
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_169
timestamp 1644511149
transform 1 0 16652 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_175
timestamp 1644511149
transform 1 0 17204 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_180
timestamp 1644511149
transform 1 0 17664 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_186
timestamp 1644511149
transform 1 0 18216 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_192
timestamp 1644511149
transform 1 0 18768 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_197
timestamp 1644511149
transform 1 0 19228 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_203
timestamp 1644511149
transform 1 0 19780 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_208
timestamp 1644511149
transform 1 0 20240 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_220
timestamp 1644511149
transform 1 0 21344 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_225
timestamp 1644511149
transform 1 0 21804 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_230
timestamp 1644511149
transform 1 0 22264 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_234
timestamp 1644511149
transform 1 0 22632 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_238
timestamp 1644511149
transform 1 0 23000 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_250
timestamp 1644511149
transform 1 0 24104 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_254
timestamp 1644511149
transform 1 0 24472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_259
timestamp 1644511149
transform 1 0 24932 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_263
timestamp 1644511149
transform 1 0 25300 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_275
timestamp 1644511149
transform 1 0 26404 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1644511149
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_281
timestamp 1644511149
transform 1 0 26956 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_287
timestamp 1644511149
transform 1 0 27508 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_291
timestamp 1644511149
transform 1 0 27876 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_303
timestamp 1644511149
transform 1 0 28980 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_309
timestamp 1644511149
transform 1 0 29532 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_314
timestamp 1644511149
transform 1 0 29992 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_318
timestamp 1644511149
transform 1 0 30360 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_326
timestamp 1644511149
transform 1 0 31096 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_330
timestamp 1644511149
transform 1 0 31464 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_334
timestamp 1644511149
transform 1 0 31832 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_337
timestamp 1644511149
transform 1 0 32108 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_343
timestamp 1644511149
transform 1 0 32660 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_350
timestamp 1644511149
transform 1 0 33304 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_362
timestamp 1644511149
transform 1 0 34408 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_7
timestamp 1644511149
transform 1 0 1748 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_13
timestamp 1644511149
transform 1 0 2300 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_18
timestamp 1644511149
transform 1 0 2760 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_22
timestamp 1644511149
transform 1 0 3128 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_31
timestamp 1644511149
transform 1 0 3956 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_35
timestamp 1644511149
transform 1 0 4324 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_47
timestamp 1644511149
transform 1 0 5428 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_59
timestamp 1644511149
transform 1 0 6532 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_71
timestamp 1644511149
transform 1 0 7636 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_75
timestamp 1644511149
transform 1 0 8004 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_78
timestamp 1644511149
transform 1 0 8280 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_2_85
timestamp 1644511149
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_97
timestamp 1644511149
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_109
timestamp 1644511149
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_121
timestamp 1644511149
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1644511149
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1644511149
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_141
timestamp 1644511149
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_153
timestamp 1644511149
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_165
timestamp 1644511149
transform 1 0 16284 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_172
timestamp 1644511149
transform 1 0 16928 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_180
timestamp 1644511149
transform 1 0 17664 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_185
timestamp 1644511149
transform 1 0 18124 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_190
timestamp 1644511149
transform 1 0 18584 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_199
timestamp 1644511149
transform 1 0 19412 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_203
timestamp 1644511149
transform 1 0 19780 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_215
timestamp 1644511149
transform 1 0 20884 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_227
timestamp 1644511149
transform 1 0 21988 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_239
timestamp 1644511149
transform 1 0 23092 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1644511149
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_253
timestamp 1644511149
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_265
timestamp 1644511149
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_277
timestamp 1644511149
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_289
timestamp 1644511149
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 1644511149
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1644511149
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_309
timestamp 1644511149
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_321
timestamp 1644511149
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_333
timestamp 1644511149
transform 1 0 31740 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_339
timestamp 1644511149
transform 1 0 32292 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_342
timestamp 1644511149
transform 1 0 32568 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_346
timestamp 1644511149
transform 1 0 32936 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_350
timestamp 1644511149
transform 1 0 33304 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_356
timestamp 1644511149
transform 1 0 33856 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_362
timestamp 1644511149
transform 1 0 34408 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_6
timestamp 1644511149
transform 1 0 1656 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_11
timestamp 1644511149
transform 1 0 2116 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1644511149
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1644511149
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1644511149
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1644511149
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1644511149
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_57
timestamp 1644511149
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_69
timestamp 1644511149
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_81
timestamp 1644511149
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_93
timestamp 1644511149
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1644511149
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1644511149
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_113
timestamp 1644511149
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_125
timestamp 1644511149
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_137
timestamp 1644511149
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_149
timestamp 1644511149
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1644511149
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1644511149
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_169
timestamp 1644511149
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_181
timestamp 1644511149
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_193
timestamp 1644511149
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_205
timestamp 1644511149
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1644511149
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1644511149
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_225
timestamp 1644511149
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_237
timestamp 1644511149
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_249
timestamp 1644511149
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_261
timestamp 1644511149
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1644511149
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1644511149
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_281
timestamp 1644511149
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_293
timestamp 1644511149
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_305
timestamp 1644511149
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_317
timestamp 1644511149
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1644511149
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1644511149
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_337
timestamp 1644511149
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_349
timestamp 1644511149
transform 1 0 33212 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_352
timestamp 1644511149
transform 1 0 33488 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_356
timestamp 1644511149
transform 1 0 33856 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_362
timestamp 1644511149
transform 1 0 34408 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_5
timestamp 1644511149
transform 1 0 1564 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_17
timestamp 1644511149
transform 1 0 2668 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_25
timestamp 1644511149
transform 1 0 3404 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_29
timestamp 1644511149
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_41
timestamp 1644511149
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_53
timestamp 1644511149
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_65
timestamp 1644511149
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1644511149
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1644511149
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_85
timestamp 1644511149
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_97
timestamp 1644511149
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_109
timestamp 1644511149
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_121
timestamp 1644511149
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1644511149
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1644511149
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_141
timestamp 1644511149
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_153
timestamp 1644511149
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_165
timestamp 1644511149
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_177
timestamp 1644511149
transform 1 0 17388 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_181
timestamp 1644511149
transform 1 0 17756 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_186
timestamp 1644511149
transform 1 0 18216 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_192
timestamp 1644511149
transform 1 0 18768 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_197
timestamp 1644511149
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_209
timestamp 1644511149
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_221
timestamp 1644511149
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_233
timestamp 1644511149
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1644511149
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1644511149
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_253
timestamp 1644511149
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_265
timestamp 1644511149
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_277
timestamp 1644511149
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_289
timestamp 1644511149
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1644511149
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1644511149
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_309
timestamp 1644511149
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_321
timestamp 1644511149
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_333
timestamp 1644511149
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_345
timestamp 1644511149
transform 1 0 32844 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_353
timestamp 1644511149
transform 1 0 33580 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_356
timestamp 1644511149
transform 1 0 33856 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_362
timestamp 1644511149
transform 1 0 34408 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_7
timestamp 1644511149
transform 1 0 1748 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_19
timestamp 1644511149
transform 1 0 2852 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_31
timestamp 1644511149
transform 1 0 3956 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_43
timestamp 1644511149
transform 1 0 5060 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1644511149
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_57
timestamp 1644511149
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_69
timestamp 1644511149
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_81
timestamp 1644511149
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_93
timestamp 1644511149
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_105
timestamp 1644511149
transform 1 0 10764 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_110
timestamp 1644511149
transform 1 0 11224 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_113
timestamp 1644511149
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_125
timestamp 1644511149
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_137
timestamp 1644511149
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_149
timestamp 1644511149
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1644511149
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1644511149
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_169
timestamp 1644511149
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_181
timestamp 1644511149
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_193
timestamp 1644511149
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_205
timestamp 1644511149
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1644511149
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1644511149
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_225
timestamp 1644511149
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_237
timestamp 1644511149
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_249
timestamp 1644511149
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_261
timestamp 1644511149
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1644511149
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1644511149
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_281
timestamp 1644511149
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_293
timestamp 1644511149
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_305
timestamp 1644511149
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_317
timestamp 1644511149
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1644511149
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1644511149
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_337
timestamp 1644511149
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_349
timestamp 1644511149
transform 1 0 33212 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_362
timestamp 1644511149
transform 1 0 34408 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1644511149
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1644511149
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1644511149
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_29
timestamp 1644511149
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_41
timestamp 1644511149
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_53
timestamp 1644511149
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_65
timestamp 1644511149
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1644511149
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1644511149
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_85
timestamp 1644511149
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_97
timestamp 1644511149
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_109
timestamp 1644511149
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_121
timestamp 1644511149
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1644511149
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1644511149
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_141
timestamp 1644511149
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_153
timestamp 1644511149
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_165
timestamp 1644511149
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_177
timestamp 1644511149
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1644511149
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1644511149
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_197
timestamp 1644511149
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_209
timestamp 1644511149
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_221
timestamp 1644511149
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_233
timestamp 1644511149
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1644511149
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1644511149
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_253
timestamp 1644511149
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_265
timestamp 1644511149
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_277
timestamp 1644511149
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_289
timestamp 1644511149
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1644511149
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1644511149
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_309
timestamp 1644511149
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_321
timestamp 1644511149
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_333
timestamp 1644511149
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_345
timestamp 1644511149
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_357
timestamp 1644511149
transform 1 0 33948 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_362
timestamp 1644511149
transform 1 0 34408 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_7
timestamp 1644511149
transform 1 0 1748 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_19
timestamp 1644511149
transform 1 0 2852 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_31
timestamp 1644511149
transform 1 0 3956 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_43
timestamp 1644511149
transform 1 0 5060 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1644511149
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_57
timestamp 1644511149
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_69
timestamp 1644511149
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_81
timestamp 1644511149
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_93
timestamp 1644511149
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1644511149
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1644511149
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_113
timestamp 1644511149
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_125
timestamp 1644511149
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_137
timestamp 1644511149
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_149
timestamp 1644511149
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1644511149
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1644511149
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_169
timestamp 1644511149
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_181
timestamp 1644511149
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_193
timestamp 1644511149
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_205
timestamp 1644511149
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1644511149
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1644511149
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_225
timestamp 1644511149
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_237
timestamp 1644511149
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_249
timestamp 1644511149
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_261
timestamp 1644511149
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1644511149
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1644511149
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_281
timestamp 1644511149
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_293
timestamp 1644511149
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_305
timestamp 1644511149
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_317
timestamp 1644511149
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1644511149
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1644511149
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_337
timestamp 1644511149
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_349
timestamp 1644511149
transform 1 0 33212 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_353
timestamp 1644511149
transform 1 0 33580 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_356
timestamp 1644511149
transform 1 0 33856 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_362
timestamp 1644511149
transform 1 0 34408 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1644511149
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1644511149
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1644511149
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_29
timestamp 1644511149
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_41
timestamp 1644511149
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_53
timestamp 1644511149
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_65
timestamp 1644511149
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1644511149
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1644511149
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_85
timestamp 1644511149
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_97
timestamp 1644511149
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_109
timestamp 1644511149
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_121
timestamp 1644511149
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1644511149
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1644511149
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_141
timestamp 1644511149
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_153
timestamp 1644511149
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_165
timestamp 1644511149
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_177
timestamp 1644511149
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1644511149
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1644511149
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_197
timestamp 1644511149
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_209
timestamp 1644511149
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_221
timestamp 1644511149
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_233
timestamp 1644511149
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1644511149
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1644511149
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_253
timestamp 1644511149
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_265
timestamp 1644511149
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_277
timestamp 1644511149
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_289
timestamp 1644511149
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1644511149
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1644511149
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_309
timestamp 1644511149
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_321
timestamp 1644511149
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_333
timestamp 1644511149
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_345
timestamp 1644511149
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1644511149
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1644511149
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_7
timestamp 1644511149
transform 1 0 1748 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_11
timestamp 1644511149
transform 1 0 2116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_23
timestamp 1644511149
transform 1 0 3220 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_35
timestamp 1644511149
transform 1 0 4324 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_47
timestamp 1644511149
transform 1 0 5428 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1644511149
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_57
timestamp 1644511149
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_69
timestamp 1644511149
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_81
timestamp 1644511149
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_93
timestamp 1644511149
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1644511149
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1644511149
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_113
timestamp 1644511149
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_125
timestamp 1644511149
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_137
timestamp 1644511149
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_149
timestamp 1644511149
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1644511149
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1644511149
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_169
timestamp 1644511149
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_181
timestamp 1644511149
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_193
timestamp 1644511149
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_205
timestamp 1644511149
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1644511149
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1644511149
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_225
timestamp 1644511149
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_237
timestamp 1644511149
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_249
timestamp 1644511149
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_261
timestamp 1644511149
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1644511149
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1644511149
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_281
timestamp 1644511149
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_293
timestamp 1644511149
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_305
timestamp 1644511149
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_317
timestamp 1644511149
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1644511149
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1644511149
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_337
timestamp 1644511149
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_349
timestamp 1644511149
transform 1 0 33212 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_357
timestamp 1644511149
transform 1 0 33948 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_362
timestamp 1644511149
transform 1 0 34408 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_7
timestamp 1644511149
transform 1 0 1748 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_19
timestamp 1644511149
transform 1 0 2852 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1644511149
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_29
timestamp 1644511149
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_41
timestamp 1644511149
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_53
timestamp 1644511149
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_65
timestamp 1644511149
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1644511149
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1644511149
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_85
timestamp 1644511149
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_97
timestamp 1644511149
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_109
timestamp 1644511149
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_121
timestamp 1644511149
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1644511149
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1644511149
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_141
timestamp 1644511149
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_153
timestamp 1644511149
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_165
timestamp 1644511149
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_177
timestamp 1644511149
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1644511149
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1644511149
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_197
timestamp 1644511149
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_209
timestamp 1644511149
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_221
timestamp 1644511149
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_233
timestamp 1644511149
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1644511149
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1644511149
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_253
timestamp 1644511149
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_265
timestamp 1644511149
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_277
timestamp 1644511149
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_289
timestamp 1644511149
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1644511149
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1644511149
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_309
timestamp 1644511149
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_321
timestamp 1644511149
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_333
timestamp 1644511149
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_345
timestamp 1644511149
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_357
timestamp 1644511149
transform 1 0 33948 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_362
timestamp 1644511149
transform 1 0 34408 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1644511149
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1644511149
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_27
timestamp 1644511149
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_39
timestamp 1644511149
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1644511149
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1644511149
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_57
timestamp 1644511149
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_69
timestamp 1644511149
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_81
timestamp 1644511149
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_93
timestamp 1644511149
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1644511149
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1644511149
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_113
timestamp 1644511149
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_125
timestamp 1644511149
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_137
timestamp 1644511149
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_149
timestamp 1644511149
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1644511149
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1644511149
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_169
timestamp 1644511149
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_181
timestamp 1644511149
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_193
timestamp 1644511149
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_205
timestamp 1644511149
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1644511149
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1644511149
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_225
timestamp 1644511149
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_237
timestamp 1644511149
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_249
timestamp 1644511149
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_261
timestamp 1644511149
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1644511149
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1644511149
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_281
timestamp 1644511149
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_293
timestamp 1644511149
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_305
timestamp 1644511149
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_317
timestamp 1644511149
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1644511149
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1644511149
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_337
timestamp 1644511149
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_349
timestamp 1644511149
transform 1 0 33212 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_353
timestamp 1644511149
transform 1 0 33580 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_356
timestamp 1644511149
transform 1 0 33856 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_362
timestamp 1644511149
transform 1 0 34408 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_7
timestamp 1644511149
transform 1 0 1748 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_11
timestamp 1644511149
transform 1 0 2116 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_23
timestamp 1644511149
transform 1 0 3220 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1644511149
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_29
timestamp 1644511149
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_41
timestamp 1644511149
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_53
timestamp 1644511149
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_65
timestamp 1644511149
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1644511149
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1644511149
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_85
timestamp 1644511149
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_97
timestamp 1644511149
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_109
timestamp 1644511149
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_121
timestamp 1644511149
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1644511149
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1644511149
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_141
timestamp 1644511149
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_153
timestamp 1644511149
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_165
timestamp 1644511149
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_177
timestamp 1644511149
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1644511149
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1644511149
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_197
timestamp 1644511149
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_209
timestamp 1644511149
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_221
timestamp 1644511149
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_233
timestamp 1644511149
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1644511149
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1644511149
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_253
timestamp 1644511149
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_265
timestamp 1644511149
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_277
timestamp 1644511149
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_289
timestamp 1644511149
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1644511149
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1644511149
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_309
timestamp 1644511149
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_321
timestamp 1644511149
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_333
timestamp 1644511149
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_345
timestamp 1644511149
transform 1 0 32844 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_353
timestamp 1644511149
transform 1 0 33580 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_356
timestamp 1644511149
transform 1 0 33856 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_362
timestamp 1644511149
transform 1 0 34408 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1644511149
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1644511149
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1644511149
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_39
timestamp 1644511149
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1644511149
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1644511149
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_57
timestamp 1644511149
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_69
timestamp 1644511149
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_81
timestamp 1644511149
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_93
timestamp 1644511149
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1644511149
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1644511149
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_113
timestamp 1644511149
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_125
timestamp 1644511149
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_137
timestamp 1644511149
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_149
timestamp 1644511149
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1644511149
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1644511149
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_169
timestamp 1644511149
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_181
timestamp 1644511149
transform 1 0 17756 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_186
timestamp 1644511149
transform 1 0 18216 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_190
timestamp 1644511149
transform 1 0 18584 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_202
timestamp 1644511149
transform 1 0 19688 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_214
timestamp 1644511149
transform 1 0 20792 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_222
timestamp 1644511149
transform 1 0 21528 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_225
timestamp 1644511149
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_237
timestamp 1644511149
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_249
timestamp 1644511149
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_261
timestamp 1644511149
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1644511149
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1644511149
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_281
timestamp 1644511149
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_293
timestamp 1644511149
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_305
timestamp 1644511149
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_317
timestamp 1644511149
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1644511149
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1644511149
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_337
timestamp 1644511149
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_349
timestamp 1644511149
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_361
timestamp 1644511149
transform 1 0 34316 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1644511149
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1644511149
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1644511149
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_29
timestamp 1644511149
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_41
timestamp 1644511149
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_53
timestamp 1644511149
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_65
timestamp 1644511149
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1644511149
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1644511149
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_85
timestamp 1644511149
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_97
timestamp 1644511149
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_109
timestamp 1644511149
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_121
timestamp 1644511149
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1644511149
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1644511149
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_141
timestamp 1644511149
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_153
timestamp 1644511149
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_165
timestamp 1644511149
transform 1 0 16284 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_173
timestamp 1644511149
transform 1 0 17020 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_180
timestamp 1644511149
transform 1 0 17664 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_192
timestamp 1644511149
transform 1 0 18768 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_197
timestamp 1644511149
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_209
timestamp 1644511149
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_221
timestamp 1644511149
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_233
timestamp 1644511149
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1644511149
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1644511149
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_253
timestamp 1644511149
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_265
timestamp 1644511149
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_277
timestamp 1644511149
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_289
timestamp 1644511149
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_301
timestamp 1644511149
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1644511149
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_309
timestamp 1644511149
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_321
timestamp 1644511149
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_333
timestamp 1644511149
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_345
timestamp 1644511149
transform 1 0 32844 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_353
timestamp 1644511149
transform 1 0 33580 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_357
timestamp 1644511149
transform 1 0 33948 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_362
timestamp 1644511149
transform 1 0 34408 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_6
timestamp 1644511149
transform 1 0 1656 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_10
timestamp 1644511149
transform 1 0 2024 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_22
timestamp 1644511149
transform 1 0 3128 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_34
timestamp 1644511149
transform 1 0 4232 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_46
timestamp 1644511149
transform 1 0 5336 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_54
timestamp 1644511149
transform 1 0 6072 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_57
timestamp 1644511149
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_69
timestamp 1644511149
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_81
timestamp 1644511149
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_93
timestamp 1644511149
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1644511149
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1644511149
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_113
timestamp 1644511149
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_125
timestamp 1644511149
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_137
timestamp 1644511149
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_149
timestamp 1644511149
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1644511149
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1644511149
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_169
timestamp 1644511149
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_181
timestamp 1644511149
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_193
timestamp 1644511149
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_205
timestamp 1644511149
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1644511149
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1644511149
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_225
timestamp 1644511149
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_237
timestamp 1644511149
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_249
timestamp 1644511149
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_261
timestamp 1644511149
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp 1644511149
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1644511149
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_281
timestamp 1644511149
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_293
timestamp 1644511149
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_305
timestamp 1644511149
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_317
timestamp 1644511149
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_329
timestamp 1644511149
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1644511149
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_337
timestamp 1644511149
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_349
timestamp 1644511149
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_361
timestamp 1644511149
transform 1 0 34316 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_5
timestamp 1644511149
transform 1 0 1564 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_17
timestamp 1644511149
transform 1 0 2668 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_25
timestamp 1644511149
transform 1 0 3404 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_29
timestamp 1644511149
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_41
timestamp 1644511149
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_53
timestamp 1644511149
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_65
timestamp 1644511149
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1644511149
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1644511149
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_85
timestamp 1644511149
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_97
timestamp 1644511149
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_109
timestamp 1644511149
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_121
timestamp 1644511149
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1644511149
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1644511149
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_141
timestamp 1644511149
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_153
timestamp 1644511149
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_165
timestamp 1644511149
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_177
timestamp 1644511149
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1644511149
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1644511149
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_197
timestamp 1644511149
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_209
timestamp 1644511149
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_221
timestamp 1644511149
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_233
timestamp 1644511149
transform 1 0 22540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_245
timestamp 1644511149
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1644511149
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_253
timestamp 1644511149
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_265
timestamp 1644511149
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_277
timestamp 1644511149
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_289
timestamp 1644511149
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_301
timestamp 1644511149
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1644511149
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_309
timestamp 1644511149
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_321
timestamp 1644511149
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_333
timestamp 1644511149
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_345
timestamp 1644511149
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_357
timestamp 1644511149
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1644511149
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_13
timestamp 1644511149
transform 1 0 2300 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_25
timestamp 1644511149
transform 1 0 3404 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_37
timestamp 1644511149
transform 1 0 4508 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_49
timestamp 1644511149
transform 1 0 5612 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1644511149
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_57
timestamp 1644511149
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_69
timestamp 1644511149
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_81
timestamp 1644511149
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_93
timestamp 1644511149
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1644511149
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1644511149
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_113
timestamp 1644511149
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_125
timestamp 1644511149
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_137
timestamp 1644511149
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_149
timestamp 1644511149
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1644511149
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1644511149
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_169
timestamp 1644511149
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_181
timestamp 1644511149
transform 1 0 17756 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_186
timestamp 1644511149
transform 1 0 18216 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_198
timestamp 1644511149
transform 1 0 19320 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_210
timestamp 1644511149
transform 1 0 20424 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_222
timestamp 1644511149
transform 1 0 21528 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_225
timestamp 1644511149
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_237
timestamp 1644511149
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_249
timestamp 1644511149
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_261
timestamp 1644511149
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 1644511149
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1644511149
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_281
timestamp 1644511149
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_293
timestamp 1644511149
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_305
timestamp 1644511149
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_317
timestamp 1644511149
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_329
timestamp 1644511149
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1644511149
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_337
timestamp 1644511149
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_349
timestamp 1644511149
transform 1 0 33212 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_357
timestamp 1644511149
transform 1 0 33948 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_362
timestamp 1644511149
transform 1 0 34408 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1644511149
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1644511149
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1644511149
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_29
timestamp 1644511149
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_41
timestamp 1644511149
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_53
timestamp 1644511149
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_65
timestamp 1644511149
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1644511149
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1644511149
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_85
timestamp 1644511149
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_97
timestamp 1644511149
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_109
timestamp 1644511149
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_121
timestamp 1644511149
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1644511149
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1644511149
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_141
timestamp 1644511149
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_153
timestamp 1644511149
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_165
timestamp 1644511149
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_177
timestamp 1644511149
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 1644511149
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1644511149
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_197
timestamp 1644511149
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_209
timestamp 1644511149
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_221
timestamp 1644511149
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_233
timestamp 1644511149
transform 1 0 22540 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_245
timestamp 1644511149
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1644511149
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_253
timestamp 1644511149
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_265
timestamp 1644511149
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_277
timestamp 1644511149
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_289
timestamp 1644511149
transform 1 0 27692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_301
timestamp 1644511149
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1644511149
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_309
timestamp 1644511149
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_321
timestamp 1644511149
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_333
timestamp 1644511149
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_345
timestamp 1644511149
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 1644511149
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1644511149
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_7
timestamp 1644511149
transform 1 0 1748 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_11
timestamp 1644511149
transform 1 0 2116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_23
timestamp 1644511149
transform 1 0 3220 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_35
timestamp 1644511149
transform 1 0 4324 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_47
timestamp 1644511149
transform 1 0 5428 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1644511149
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_57
timestamp 1644511149
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_69
timestamp 1644511149
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_81
timestamp 1644511149
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_93
timestamp 1644511149
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1644511149
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1644511149
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_113
timestamp 1644511149
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_125
timestamp 1644511149
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_137
timestamp 1644511149
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_149
timestamp 1644511149
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1644511149
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1644511149
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_169
timestamp 1644511149
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_181
timestamp 1644511149
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_193
timestamp 1644511149
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_205
timestamp 1644511149
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_217
timestamp 1644511149
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1644511149
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_225
timestamp 1644511149
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_237
timestamp 1644511149
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_249
timestamp 1644511149
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_261
timestamp 1644511149
transform 1 0 25116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_273
timestamp 1644511149
transform 1 0 26220 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1644511149
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_281
timestamp 1644511149
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_293
timestamp 1644511149
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_305
timestamp 1644511149
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_317
timestamp 1644511149
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_329
timestamp 1644511149
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1644511149
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_337
timestamp 1644511149
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_349
timestamp 1644511149
transform 1 0 33212 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_353
timestamp 1644511149
transform 1 0 33580 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_356
timestamp 1644511149
transform 1 0 33856 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_362
timestamp 1644511149
transform 1 0 34408 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1644511149
transform 1 0 1380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_9
timestamp 1644511149
transform 1 0 1932 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_13
timestamp 1644511149
transform 1 0 2300 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_25
timestamp 1644511149
transform 1 0 3404 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_29
timestamp 1644511149
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_41
timestamp 1644511149
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_53
timestamp 1644511149
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_65
timestamp 1644511149
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1644511149
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1644511149
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_85
timestamp 1644511149
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_97
timestamp 1644511149
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_109
timestamp 1644511149
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_121
timestamp 1644511149
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1644511149
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1644511149
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_141
timestamp 1644511149
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_153
timestamp 1644511149
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_165
timestamp 1644511149
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_177
timestamp 1644511149
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_189
timestamp 1644511149
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1644511149
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_197
timestamp 1644511149
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_209
timestamp 1644511149
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_221
timestamp 1644511149
transform 1 0 21436 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_233
timestamp 1644511149
transform 1 0 22540 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_245
timestamp 1644511149
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1644511149
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_253
timestamp 1644511149
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_265
timestamp 1644511149
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_277
timestamp 1644511149
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_289
timestamp 1644511149
transform 1 0 27692 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_301
timestamp 1644511149
transform 1 0 28796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1644511149
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_309
timestamp 1644511149
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_321
timestamp 1644511149
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_333
timestamp 1644511149
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_345
timestamp 1644511149
transform 1 0 32844 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_353
timestamp 1644511149
transform 1 0 33580 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_356
timestamp 1644511149
transform 1 0 33856 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_362
timestamp 1644511149
transform 1 0 34408 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1644511149
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1644511149
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 1644511149
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_39
timestamp 1644511149
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1644511149
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1644511149
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_57
timestamp 1644511149
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_69
timestamp 1644511149
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_81
timestamp 1644511149
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_93
timestamp 1644511149
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1644511149
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1644511149
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_113
timestamp 1644511149
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_125
timestamp 1644511149
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_137
timestamp 1644511149
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_149
timestamp 1644511149
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 1644511149
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1644511149
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_169
timestamp 1644511149
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_181
timestamp 1644511149
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_193
timestamp 1644511149
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_205
timestamp 1644511149
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_217
timestamp 1644511149
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1644511149
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_225
timestamp 1644511149
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_237
timestamp 1644511149
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_249
timestamp 1644511149
transform 1 0 24012 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_261
timestamp 1644511149
transform 1 0 25116 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_273
timestamp 1644511149
transform 1 0 26220 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1644511149
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_281
timestamp 1644511149
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_293
timestamp 1644511149
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_305
timestamp 1644511149
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_317
timestamp 1644511149
transform 1 0 30268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_329
timestamp 1644511149
transform 1 0 31372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1644511149
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_337
timestamp 1644511149
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_349
timestamp 1644511149
transform 1 0 33212 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_362
timestamp 1644511149
transform 1 0 34408 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_7
timestamp 1644511149
transform 1 0 1748 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_19
timestamp 1644511149
transform 1 0 2852 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1644511149
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_29
timestamp 1644511149
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_41
timestamp 1644511149
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_53
timestamp 1644511149
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_65
timestamp 1644511149
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1644511149
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1644511149
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_85
timestamp 1644511149
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_97
timestamp 1644511149
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_109
timestamp 1644511149
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_121
timestamp 1644511149
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1644511149
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1644511149
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_141
timestamp 1644511149
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_153
timestamp 1644511149
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_165
timestamp 1644511149
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_177
timestamp 1644511149
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_189
timestamp 1644511149
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1644511149
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_197
timestamp 1644511149
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_209
timestamp 1644511149
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_221
timestamp 1644511149
transform 1 0 21436 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_233
timestamp 1644511149
transform 1 0 22540 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_245
timestamp 1644511149
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1644511149
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_253
timestamp 1644511149
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_265
timestamp 1644511149
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_277
timestamp 1644511149
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_289
timestamp 1644511149
transform 1 0 27692 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_301
timestamp 1644511149
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1644511149
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_309
timestamp 1644511149
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_321
timestamp 1644511149
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_333
timestamp 1644511149
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_345
timestamp 1644511149
transform 1 0 32844 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_22_353
timestamp 1644511149
transform 1 0 33580 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_357
timestamp 1644511149
transform 1 0 33948 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_362
timestamp 1644511149
transform 1 0 34408 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1644511149
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1644511149
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_27
timestamp 1644511149
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_39
timestamp 1644511149
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1644511149
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1644511149
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_57
timestamp 1644511149
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_69
timestamp 1644511149
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_81
timestamp 1644511149
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_93
timestamp 1644511149
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1644511149
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1644511149
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_113
timestamp 1644511149
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_125
timestamp 1644511149
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_137
timestamp 1644511149
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_149
timestamp 1644511149
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1644511149
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1644511149
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_169
timestamp 1644511149
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_181
timestamp 1644511149
transform 1 0 17756 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_186
timestamp 1644511149
transform 1 0 18216 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_192
timestamp 1644511149
transform 1 0 18768 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_196
timestamp 1644511149
transform 1 0 19136 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_208
timestamp 1644511149
transform 1 0 20240 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_220
timestamp 1644511149
transform 1 0 21344 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_225
timestamp 1644511149
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_237
timestamp 1644511149
transform 1 0 22908 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_249
timestamp 1644511149
transform 1 0 24012 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_261
timestamp 1644511149
transform 1 0 25116 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_273
timestamp 1644511149
transform 1 0 26220 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 1644511149
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_281
timestamp 1644511149
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_293
timestamp 1644511149
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_305
timestamp 1644511149
transform 1 0 29164 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_317
timestamp 1644511149
transform 1 0 30268 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_329
timestamp 1644511149
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1644511149
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_337
timestamp 1644511149
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_349
timestamp 1644511149
transform 1 0 33212 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_360
timestamp 1644511149
transform 1 0 34224 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_6
timestamp 1644511149
transform 1 0 1656 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_10
timestamp 1644511149
transform 1 0 2024 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_22
timestamp 1644511149
transform 1 0 3128 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_24_29
timestamp 1644511149
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_41
timestamp 1644511149
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_53
timestamp 1644511149
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_65
timestamp 1644511149
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1644511149
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1644511149
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_85
timestamp 1644511149
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_97
timestamp 1644511149
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_109
timestamp 1644511149
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_121
timestamp 1644511149
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1644511149
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1644511149
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_141
timestamp 1644511149
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_153
timestamp 1644511149
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_165
timestamp 1644511149
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_177
timestamp 1644511149
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_189
timestamp 1644511149
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1644511149
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_197
timestamp 1644511149
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_209
timestamp 1644511149
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_221
timestamp 1644511149
transform 1 0 21436 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_233
timestamp 1644511149
transform 1 0 22540 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_245
timestamp 1644511149
transform 1 0 23644 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1644511149
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_253
timestamp 1644511149
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_265
timestamp 1644511149
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_277
timestamp 1644511149
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_289
timestamp 1644511149
transform 1 0 27692 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_301
timestamp 1644511149
transform 1 0 28796 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1644511149
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_309
timestamp 1644511149
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_321
timestamp 1644511149
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_333
timestamp 1644511149
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_345
timestamp 1644511149
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_357
timestamp 1644511149
transform 1 0 33948 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_362
timestamp 1644511149
transform 1 0 34408 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_7
timestamp 1644511149
transform 1 0 1748 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_19
timestamp 1644511149
transform 1 0 2852 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_31
timestamp 1644511149
transform 1 0 3956 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_43
timestamp 1644511149
transform 1 0 5060 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1644511149
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_57
timestamp 1644511149
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_69
timestamp 1644511149
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_81
timestamp 1644511149
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_93
timestamp 1644511149
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1644511149
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1644511149
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_113
timestamp 1644511149
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_125
timestamp 1644511149
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_137
timestamp 1644511149
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_149
timestamp 1644511149
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1644511149
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1644511149
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_169
timestamp 1644511149
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_181
timestamp 1644511149
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_193
timestamp 1644511149
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_205
timestamp 1644511149
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_217
timestamp 1644511149
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1644511149
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_225
timestamp 1644511149
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_237
timestamp 1644511149
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_249
timestamp 1644511149
transform 1 0 24012 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_261
timestamp 1644511149
transform 1 0 25116 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_273
timestamp 1644511149
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1644511149
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_281
timestamp 1644511149
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_293
timestamp 1644511149
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_305
timestamp 1644511149
transform 1 0 29164 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_317
timestamp 1644511149
transform 1 0 30268 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_329
timestamp 1644511149
transform 1 0 31372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1644511149
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_337
timestamp 1644511149
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_349
timestamp 1644511149
transform 1 0 33212 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_362
timestamp 1644511149
transform 1 0 34408 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1644511149
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1644511149
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1644511149
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_29
timestamp 1644511149
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_41
timestamp 1644511149
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_53
timestamp 1644511149
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_65
timestamp 1644511149
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1644511149
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1644511149
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_85
timestamp 1644511149
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_97
timestamp 1644511149
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_109
timestamp 1644511149
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_121
timestamp 1644511149
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1644511149
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1644511149
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_141
timestamp 1644511149
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_153
timestamp 1644511149
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_165
timestamp 1644511149
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_177
timestamp 1644511149
transform 1 0 17388 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_181
timestamp 1644511149
transform 1 0 17756 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_193
timestamp 1644511149
transform 1 0 18860 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_197
timestamp 1644511149
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_209
timestamp 1644511149
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_221
timestamp 1644511149
transform 1 0 21436 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_233
timestamp 1644511149
transform 1 0 22540 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_245
timestamp 1644511149
transform 1 0 23644 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1644511149
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_253
timestamp 1644511149
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_265
timestamp 1644511149
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_277
timestamp 1644511149
transform 1 0 26588 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_289
timestamp 1644511149
transform 1 0 27692 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_301
timestamp 1644511149
transform 1 0 28796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1644511149
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_309
timestamp 1644511149
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_321
timestamp 1644511149
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_333
timestamp 1644511149
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_345
timestamp 1644511149
transform 1 0 32844 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_357
timestamp 1644511149
transform 1 0 33948 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_362
timestamp 1644511149
transform 1 0 34408 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_7
timestamp 1644511149
transform 1 0 1748 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_19
timestamp 1644511149
transform 1 0 2852 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_31
timestamp 1644511149
transform 1 0 3956 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_43
timestamp 1644511149
transform 1 0 5060 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1644511149
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_57
timestamp 1644511149
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_69
timestamp 1644511149
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_81
timestamp 1644511149
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_93
timestamp 1644511149
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1644511149
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1644511149
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_113
timestamp 1644511149
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_125
timestamp 1644511149
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_137
timestamp 1644511149
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_149
timestamp 1644511149
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1644511149
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1644511149
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_169
timestamp 1644511149
transform 1 0 16652 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_179
timestamp 1644511149
transform 1 0 17572 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_185
timestamp 1644511149
transform 1 0 18124 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_191
timestamp 1644511149
transform 1 0 18676 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_195
timestamp 1644511149
transform 1 0 19044 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_207
timestamp 1644511149
transform 1 0 20148 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_219
timestamp 1644511149
transform 1 0 21252 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1644511149
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_225
timestamp 1644511149
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_237
timestamp 1644511149
transform 1 0 22908 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_249
timestamp 1644511149
transform 1 0 24012 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_261
timestamp 1644511149
transform 1 0 25116 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_273
timestamp 1644511149
transform 1 0 26220 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1644511149
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_281
timestamp 1644511149
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_293
timestamp 1644511149
transform 1 0 28060 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_305
timestamp 1644511149
transform 1 0 29164 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_311
timestamp 1644511149
transform 1 0 29716 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_315
timestamp 1644511149
transform 1 0 30084 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_327
timestamp 1644511149
transform 1 0 31188 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 1644511149
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_337
timestamp 1644511149
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_349
timestamp 1644511149
transform 1 0 33212 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_356
timestamp 1644511149
transform 1 0 33856 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_362
timestamp 1644511149
transform 1 0 34408 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_3
timestamp 1644511149
transform 1 0 1380 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_10
timestamp 1644511149
transform 1 0 2024 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_18
timestamp 1644511149
transform 1 0 2760 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_26
timestamp 1644511149
transform 1 0 3496 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_29
timestamp 1644511149
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_41
timestamp 1644511149
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_53
timestamp 1644511149
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_65
timestamp 1644511149
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1644511149
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1644511149
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_85
timestamp 1644511149
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_97
timestamp 1644511149
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_109
timestamp 1644511149
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_121
timestamp 1644511149
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1644511149
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1644511149
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_141
timestamp 1644511149
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_153
timestamp 1644511149
transform 1 0 15180 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_161
timestamp 1644511149
transform 1 0 15916 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_164
timestamp 1644511149
transform 1 0 16192 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_170
timestamp 1644511149
transform 1 0 16744 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_174
timestamp 1644511149
transform 1 0 17112 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_180
timestamp 1644511149
transform 1 0 17664 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_186
timestamp 1644511149
transform 1 0 18216 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_192
timestamp 1644511149
transform 1 0 18768 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_197
timestamp 1644511149
transform 1 0 19228 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_203
timestamp 1644511149
transform 1 0 19780 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_215
timestamp 1644511149
transform 1 0 20884 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_227
timestamp 1644511149
transform 1 0 21988 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_239
timestamp 1644511149
transform 1 0 23092 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1644511149
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_253
timestamp 1644511149
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_265
timestamp 1644511149
transform 1 0 25484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_277
timestamp 1644511149
transform 1 0 26588 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_289
timestamp 1644511149
transform 1 0 27692 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_301
timestamp 1644511149
transform 1 0 28796 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp 1644511149
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_309
timestamp 1644511149
transform 1 0 29532 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_315
timestamp 1644511149
transform 1 0 30084 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_319
timestamp 1644511149
transform 1 0 30452 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_331
timestamp 1644511149
transform 1 0 31556 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_343
timestamp 1644511149
transform 1 0 32660 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_355
timestamp 1644511149
transform 1 0 33764 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1644511149
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_3
timestamp 1644511149
transform 1 0 1380 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_10
timestamp 1644511149
transform 1 0 2024 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_15
timestamp 1644511149
transform 1 0 2484 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_23
timestamp 1644511149
transform 1 0 3220 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_29
timestamp 1644511149
transform 1 0 3772 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_41
timestamp 1644511149
transform 1 0 4876 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 1644511149
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1644511149
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_57
timestamp 1644511149
transform 1 0 6348 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_63
timestamp 1644511149
transform 1 0 6900 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_68
timestamp 1644511149
transform 1 0 7360 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_80
timestamp 1644511149
transform 1 0 8464 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_92
timestamp 1644511149
transform 1 0 9568 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_104
timestamp 1644511149
transform 1 0 10672 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_29_113
timestamp 1644511149
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_125
timestamp 1644511149
transform 1 0 12604 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_131
timestamp 1644511149
transform 1 0 13156 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_143
timestamp 1644511149
transform 1 0 14260 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_155
timestamp 1644511149
transform 1 0 15364 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_162
timestamp 1644511149
transform 1 0 16008 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_166
timestamp 1644511149
transform 1 0 16376 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_173
timestamp 1644511149
transform 1 0 17020 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_179
timestamp 1644511149
transform 1 0 17572 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_185
timestamp 1644511149
transform 1 0 18124 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_191
timestamp 1644511149
transform 1 0 18676 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_197
timestamp 1644511149
transform 1 0 19228 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_203
timestamp 1644511149
transform 1 0 19780 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_207
timestamp 1644511149
transform 1 0 20148 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_219
timestamp 1644511149
transform 1 0 21252 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1644511149
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_225
timestamp 1644511149
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_237
timestamp 1644511149
transform 1 0 22908 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_249
timestamp 1644511149
transform 1 0 24012 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_257
timestamp 1644511149
transform 1 0 24748 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_269
timestamp 1644511149
transform 1 0 25852 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_277
timestamp 1644511149
transform 1 0 26588 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_281
timestamp 1644511149
transform 1 0 26956 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_289
timestamp 1644511149
transform 1 0 27692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_301
timestamp 1644511149
transform 1 0 28796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_310
timestamp 1644511149
transform 1 0 29624 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_316
timestamp 1644511149
transform 1 0 30176 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_320
timestamp 1644511149
transform 1 0 30544 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_29_330
timestamp 1644511149
transform 1 0 31464 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_29_337
timestamp 1644511149
transform 1 0 32108 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_343
timestamp 1644511149
transform 1 0 32660 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_351
timestamp 1644511149
transform 1 0 33396 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_356
timestamp 1644511149
transform 1 0 33856 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_362
timestamp 1644511149
transform 1 0 34408 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_7
timestamp 1644511149
transform 1 0 1748 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_12
timestamp 1644511149
transform 1 0 2208 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_16
timestamp 1644511149
transform 1 0 2576 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_29
timestamp 1644511149
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_41
timestamp 1644511149
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_53
timestamp 1644511149
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_65
timestamp 1644511149
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1644511149
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1644511149
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_85
timestamp 1644511149
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_97
timestamp 1644511149
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_109
timestamp 1644511149
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_121
timestamp 1644511149
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1644511149
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1644511149
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_141
timestamp 1644511149
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_153
timestamp 1644511149
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_165
timestamp 1644511149
transform 1 0 16284 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_171
timestamp 1644511149
transform 1 0 16836 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_174
timestamp 1644511149
transform 1 0 17112 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_180
timestamp 1644511149
transform 1 0 17664 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_186
timestamp 1644511149
transform 1 0 18216 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_192
timestamp 1644511149
transform 1 0 18768 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_199
timestamp 1644511149
transform 1 0 19412 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_211
timestamp 1644511149
transform 1 0 20516 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_216
timestamp 1644511149
transform 1 0 20976 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_220
timestamp 1644511149
transform 1 0 21344 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_232
timestamp 1644511149
transform 1 0 22448 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_30_244
timestamp 1644511149
transform 1 0 23552 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_253
timestamp 1644511149
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_265
timestamp 1644511149
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_277
timestamp 1644511149
transform 1 0 26588 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_289
timestamp 1644511149
transform 1 0 27692 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_301
timestamp 1644511149
transform 1 0 28796 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_307
timestamp 1644511149
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_313
timestamp 1644511149
transform 1 0 29900 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_325
timestamp 1644511149
transform 1 0 31004 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_337
timestamp 1644511149
transform 1 0 32108 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_349
timestamp 1644511149
transform 1 0 33212 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_30_357
timestamp 1644511149
transform 1 0 33948 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_362
timestamp 1644511149
transform 1 0 34408 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_7
timestamp 1644511149
transform 1 0 1748 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_11
timestamp 1644511149
transform 1 0 2116 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_23
timestamp 1644511149
transform 1 0 3220 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_35
timestamp 1644511149
transform 1 0 4324 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_47
timestamp 1644511149
transform 1 0 5428 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1644511149
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_57
timestamp 1644511149
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_69
timestamp 1644511149
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_81
timestamp 1644511149
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_93
timestamp 1644511149
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1644511149
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1644511149
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_113
timestamp 1644511149
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_125
timestamp 1644511149
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_137
timestamp 1644511149
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_149
timestamp 1644511149
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 1644511149
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1644511149
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_169
timestamp 1644511149
transform 1 0 16652 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_173
timestamp 1644511149
transform 1 0 17020 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_176
timestamp 1644511149
transform 1 0 17296 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_186
timestamp 1644511149
transform 1 0 18216 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_192
timestamp 1644511149
transform 1 0 18768 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_196
timestamp 1644511149
transform 1 0 19136 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_208
timestamp 1644511149
transform 1 0 20240 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_220
timestamp 1644511149
transform 1 0 21344 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_225
timestamp 1644511149
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_237
timestamp 1644511149
transform 1 0 22908 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_249
timestamp 1644511149
transform 1 0 24012 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_261
timestamp 1644511149
transform 1 0 25116 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_273
timestamp 1644511149
transform 1 0 26220 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 1644511149
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_281
timestamp 1644511149
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_293
timestamp 1644511149
transform 1 0 28060 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_305
timestamp 1644511149
transform 1 0 29164 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_317
timestamp 1644511149
transform 1 0 30268 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_329
timestamp 1644511149
transform 1 0 31372 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_335
timestamp 1644511149
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_337
timestamp 1644511149
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_349
timestamp 1644511149
transform 1 0 33212 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_357
timestamp 1644511149
transform 1 0 33948 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_362
timestamp 1644511149
transform 1 0 34408 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_13
timestamp 1644511149
transform 1 0 2300 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_25
timestamp 1644511149
transform 1 0 3404 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_29
timestamp 1644511149
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_41
timestamp 1644511149
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_53
timestamp 1644511149
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_65
timestamp 1644511149
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1644511149
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1644511149
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_85
timestamp 1644511149
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_97
timestamp 1644511149
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_109
timestamp 1644511149
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_121
timestamp 1644511149
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_133
timestamp 1644511149
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1644511149
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_141
timestamp 1644511149
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_153
timestamp 1644511149
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_165
timestamp 1644511149
transform 1 0 16284 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_177
timestamp 1644511149
transform 1 0 17388 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_189
timestamp 1644511149
transform 1 0 18492 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1644511149
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_197
timestamp 1644511149
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_209
timestamp 1644511149
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_221
timestamp 1644511149
transform 1 0 21436 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_233
timestamp 1644511149
transform 1 0 22540 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_245
timestamp 1644511149
transform 1 0 23644 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1644511149
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_253
timestamp 1644511149
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_265
timestamp 1644511149
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_277
timestamp 1644511149
transform 1 0 26588 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_289
timestamp 1644511149
transform 1 0 27692 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_301
timestamp 1644511149
transform 1 0 28796 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_307
timestamp 1644511149
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_309
timestamp 1644511149
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_321
timestamp 1644511149
transform 1 0 30636 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_333
timestamp 1644511149
transform 1 0 31740 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_345
timestamp 1644511149
transform 1 0 32844 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_353
timestamp 1644511149
transform 1 0 33580 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_357
timestamp 1644511149
transform 1 0 33948 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_362
timestamp 1644511149
transform 1 0 34408 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_5
timestamp 1644511149
transform 1 0 1564 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_17
timestamp 1644511149
transform 1 0 2668 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_29
timestamp 1644511149
transform 1 0 3772 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_41
timestamp 1644511149
transform 1 0 4876 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_53
timestamp 1644511149
transform 1 0 5980 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_57
timestamp 1644511149
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_69
timestamp 1644511149
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_81
timestamp 1644511149
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_93
timestamp 1644511149
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1644511149
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1644511149
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_113
timestamp 1644511149
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_125
timestamp 1644511149
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_137
timestamp 1644511149
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_149
timestamp 1644511149
transform 1 0 14812 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_161
timestamp 1644511149
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1644511149
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_169
timestamp 1644511149
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_181
timestamp 1644511149
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_193
timestamp 1644511149
transform 1 0 18860 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_205
timestamp 1644511149
transform 1 0 19964 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_217
timestamp 1644511149
transform 1 0 21068 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1644511149
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_225
timestamp 1644511149
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_237
timestamp 1644511149
transform 1 0 22908 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_249
timestamp 1644511149
transform 1 0 24012 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_261
timestamp 1644511149
transform 1 0 25116 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_273
timestamp 1644511149
transform 1 0 26220 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1644511149
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_281
timestamp 1644511149
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_293
timestamp 1644511149
transform 1 0 28060 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_305
timestamp 1644511149
transform 1 0 29164 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_317
timestamp 1644511149
transform 1 0 30268 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_329
timestamp 1644511149
transform 1 0 31372 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_335
timestamp 1644511149
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_337
timestamp 1644511149
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_349
timestamp 1644511149
transform 1 0 33212 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_360
timestamp 1644511149
transform 1 0 34224 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1644511149
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1644511149
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1644511149
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_29
timestamp 1644511149
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_41
timestamp 1644511149
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_53
timestamp 1644511149
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_65
timestamp 1644511149
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1644511149
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1644511149
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_85
timestamp 1644511149
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_97
timestamp 1644511149
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_109
timestamp 1644511149
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_121
timestamp 1644511149
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 1644511149
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1644511149
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_141
timestamp 1644511149
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_153
timestamp 1644511149
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_165
timestamp 1644511149
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_177
timestamp 1644511149
transform 1 0 17388 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_185
timestamp 1644511149
transform 1 0 18124 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_193
timestamp 1644511149
transform 1 0 18860 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_34_197
timestamp 1644511149
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_209
timestamp 1644511149
transform 1 0 20332 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_221
timestamp 1644511149
transform 1 0 21436 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_233
timestamp 1644511149
transform 1 0 22540 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_245
timestamp 1644511149
transform 1 0 23644 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1644511149
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_253
timestamp 1644511149
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_265
timestamp 1644511149
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_277
timestamp 1644511149
transform 1 0 26588 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_289
timestamp 1644511149
transform 1 0 27692 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_301
timestamp 1644511149
transform 1 0 28796 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_307
timestamp 1644511149
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_309
timestamp 1644511149
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_321
timestamp 1644511149
transform 1 0 30636 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_333
timestamp 1644511149
transform 1 0 31740 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_345
timestamp 1644511149
transform 1 0 32844 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_350
timestamp 1644511149
transform 1 0 33304 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_362
timestamp 1644511149
transform 1 0 34408 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_7
timestamp 1644511149
transform 1 0 1748 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_19
timestamp 1644511149
transform 1 0 2852 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_31
timestamp 1644511149
transform 1 0 3956 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_43
timestamp 1644511149
transform 1 0 5060 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1644511149
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_57
timestamp 1644511149
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_69
timestamp 1644511149
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_81
timestamp 1644511149
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_93
timestamp 1644511149
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1644511149
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1644511149
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_113
timestamp 1644511149
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_125
timestamp 1644511149
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_137
timestamp 1644511149
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_149
timestamp 1644511149
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp 1644511149
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1644511149
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_169
timestamp 1644511149
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_181
timestamp 1644511149
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_193
timestamp 1644511149
transform 1 0 18860 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_205
timestamp 1644511149
transform 1 0 19964 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_217
timestamp 1644511149
transform 1 0 21068 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1644511149
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_225
timestamp 1644511149
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_237
timestamp 1644511149
transform 1 0 22908 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_249
timestamp 1644511149
transform 1 0 24012 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_261
timestamp 1644511149
transform 1 0 25116 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_273
timestamp 1644511149
transform 1 0 26220 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1644511149
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_281
timestamp 1644511149
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_293
timestamp 1644511149
transform 1 0 28060 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_305
timestamp 1644511149
transform 1 0 29164 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_317
timestamp 1644511149
transform 1 0 30268 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_329
timestamp 1644511149
transform 1 0 31372 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1644511149
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_337
timestamp 1644511149
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_349
timestamp 1644511149
transform 1 0 33212 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_362
timestamp 1644511149
transform 1 0 34408 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_3
timestamp 1644511149
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_15
timestamp 1644511149
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1644511149
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_29
timestamp 1644511149
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_41
timestamp 1644511149
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_53
timestamp 1644511149
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_65
timestamp 1644511149
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1644511149
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1644511149
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_85
timestamp 1644511149
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_97
timestamp 1644511149
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_109
timestamp 1644511149
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_121
timestamp 1644511149
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 1644511149
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1644511149
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_141
timestamp 1644511149
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_153
timestamp 1644511149
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_165
timestamp 1644511149
transform 1 0 16284 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_177
timestamp 1644511149
transform 1 0 17388 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_189
timestamp 1644511149
transform 1 0 18492 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1644511149
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_197
timestamp 1644511149
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_209
timestamp 1644511149
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_221
timestamp 1644511149
transform 1 0 21436 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_233
timestamp 1644511149
transform 1 0 22540 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_245
timestamp 1644511149
transform 1 0 23644 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1644511149
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_253
timestamp 1644511149
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_265
timestamp 1644511149
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_277
timestamp 1644511149
transform 1 0 26588 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_289
timestamp 1644511149
transform 1 0 27692 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_301
timestamp 1644511149
transform 1 0 28796 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1644511149
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_309
timestamp 1644511149
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_321
timestamp 1644511149
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_333
timestamp 1644511149
transform 1 0 31740 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_345
timestamp 1644511149
transform 1 0 32844 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_353
timestamp 1644511149
transform 1 0 33580 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_358
timestamp 1644511149
transform 1 0 34040 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_362
timestamp 1644511149
transform 1 0 34408 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_7
timestamp 1644511149
transform 1 0 1748 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_19
timestamp 1644511149
transform 1 0 2852 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_31
timestamp 1644511149
transform 1 0 3956 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_43
timestamp 1644511149
transform 1 0 5060 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1644511149
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_57
timestamp 1644511149
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_69
timestamp 1644511149
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_81
timestamp 1644511149
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_93
timestamp 1644511149
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1644511149
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1644511149
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_113
timestamp 1644511149
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_125
timestamp 1644511149
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_137
timestamp 1644511149
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_149
timestamp 1644511149
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 1644511149
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1644511149
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_169
timestamp 1644511149
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_181
timestamp 1644511149
transform 1 0 17756 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_186
timestamp 1644511149
transform 1 0 18216 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_198
timestamp 1644511149
transform 1 0 19320 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_210
timestamp 1644511149
transform 1 0 20424 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_222
timestamp 1644511149
transform 1 0 21528 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_225
timestamp 1644511149
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_237
timestamp 1644511149
transform 1 0 22908 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_249
timestamp 1644511149
transform 1 0 24012 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_261
timestamp 1644511149
transform 1 0 25116 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_273
timestamp 1644511149
transform 1 0 26220 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1644511149
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_281
timestamp 1644511149
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_293
timestamp 1644511149
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_305
timestamp 1644511149
transform 1 0 29164 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_317
timestamp 1644511149
transform 1 0 30268 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_329
timestamp 1644511149
transform 1 0 31372 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1644511149
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_337
timestamp 1644511149
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_349
timestamp 1644511149
transform 1 0 33212 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_362
timestamp 1644511149
transform 1 0 34408 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_38_3
timestamp 1644511149
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_15
timestamp 1644511149
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1644511149
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_29
timestamp 1644511149
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_41
timestamp 1644511149
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_53
timestamp 1644511149
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_65
timestamp 1644511149
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1644511149
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1644511149
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_85
timestamp 1644511149
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_97
timestamp 1644511149
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_109
timestamp 1644511149
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_121
timestamp 1644511149
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp 1644511149
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1644511149
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_141
timestamp 1644511149
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_153
timestamp 1644511149
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_165
timestamp 1644511149
transform 1 0 16284 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_177
timestamp 1644511149
transform 1 0 17388 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_189
timestamp 1644511149
transform 1 0 18492 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1644511149
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_197
timestamp 1644511149
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_209
timestamp 1644511149
transform 1 0 20332 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_221
timestamp 1644511149
transform 1 0 21436 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_233
timestamp 1644511149
transform 1 0 22540 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_245
timestamp 1644511149
transform 1 0 23644 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp 1644511149
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_253
timestamp 1644511149
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_265
timestamp 1644511149
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_277
timestamp 1644511149
transform 1 0 26588 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_289
timestamp 1644511149
transform 1 0 27692 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_301
timestamp 1644511149
transform 1 0 28796 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 1644511149
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_309
timestamp 1644511149
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_321
timestamp 1644511149
transform 1 0 30636 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_333
timestamp 1644511149
transform 1 0 31740 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_345
timestamp 1644511149
transform 1 0 32844 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_353
timestamp 1644511149
transform 1 0 33580 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_356
timestamp 1644511149
transform 1 0 33856 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_362
timestamp 1644511149
transform 1 0 34408 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_7
timestamp 1644511149
transform 1 0 1748 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_19
timestamp 1644511149
transform 1 0 2852 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_31
timestamp 1644511149
transform 1 0 3956 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_43
timestamp 1644511149
transform 1 0 5060 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1644511149
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_57
timestamp 1644511149
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_69
timestamp 1644511149
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_81
timestamp 1644511149
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_93
timestamp 1644511149
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1644511149
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1644511149
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_113
timestamp 1644511149
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_125
timestamp 1644511149
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_137
timestamp 1644511149
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_149
timestamp 1644511149
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp 1644511149
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1644511149
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_169
timestamp 1644511149
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_181
timestamp 1644511149
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_193
timestamp 1644511149
transform 1 0 18860 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_205
timestamp 1644511149
transform 1 0 19964 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_217
timestamp 1644511149
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1644511149
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_225
timestamp 1644511149
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_237
timestamp 1644511149
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_249
timestamp 1644511149
transform 1 0 24012 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_261
timestamp 1644511149
transform 1 0 25116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_273
timestamp 1644511149
transform 1 0 26220 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1644511149
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_281
timestamp 1644511149
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_293
timestamp 1644511149
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_305
timestamp 1644511149
transform 1 0 29164 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_317
timestamp 1644511149
transform 1 0 30268 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_329
timestamp 1644511149
transform 1 0 31372 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_335
timestamp 1644511149
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_337
timestamp 1644511149
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_349
timestamp 1644511149
transform 1 0 33212 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_353
timestamp 1644511149
transform 1 0 33580 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_356
timestamp 1644511149
transform 1 0 33856 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_362
timestamp 1644511149
transform 1 0 34408 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_7
timestamp 1644511149
transform 1 0 1748 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_40_11
timestamp 1644511149
transform 1 0 2116 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_23
timestamp 1644511149
transform 1 0 3220 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1644511149
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_29
timestamp 1644511149
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_41
timestamp 1644511149
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_53
timestamp 1644511149
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_65
timestamp 1644511149
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1644511149
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1644511149
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_85
timestamp 1644511149
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_97
timestamp 1644511149
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_109
timestamp 1644511149
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_121
timestamp 1644511149
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 1644511149
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1644511149
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_141
timestamp 1644511149
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_153
timestamp 1644511149
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_165
timestamp 1644511149
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_177
timestamp 1644511149
transform 1 0 17388 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_189
timestamp 1644511149
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1644511149
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_197
timestamp 1644511149
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_209
timestamp 1644511149
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_221
timestamp 1644511149
transform 1 0 21436 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_233
timestamp 1644511149
transform 1 0 22540 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_245
timestamp 1644511149
transform 1 0 23644 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1644511149
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_253
timestamp 1644511149
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_265
timestamp 1644511149
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_277
timestamp 1644511149
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_289
timestamp 1644511149
transform 1 0 27692 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_301
timestamp 1644511149
transform 1 0 28796 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 1644511149
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_309
timestamp 1644511149
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_321
timestamp 1644511149
transform 1 0 30636 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_333
timestamp 1644511149
transform 1 0 31740 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_345
timestamp 1644511149
transform 1 0 32844 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_355
timestamp 1644511149
transform 1 0 33764 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_361
timestamp 1644511149
transform 1 0 34316 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_41_7
timestamp 1644511149
transform 1 0 1748 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_11
timestamp 1644511149
transform 1 0 2116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_23
timestamp 1644511149
transform 1 0 3220 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_35
timestamp 1644511149
transform 1 0 4324 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_47
timestamp 1644511149
transform 1 0 5428 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1644511149
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_57
timestamp 1644511149
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_69
timestamp 1644511149
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_81
timestamp 1644511149
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_93
timestamp 1644511149
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1644511149
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1644511149
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_113
timestamp 1644511149
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_125
timestamp 1644511149
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_137
timestamp 1644511149
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_149
timestamp 1644511149
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_161
timestamp 1644511149
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1644511149
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_169
timestamp 1644511149
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_181
timestamp 1644511149
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_193
timestamp 1644511149
transform 1 0 18860 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_201
timestamp 1644511149
transform 1 0 19596 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_204
timestamp 1644511149
transform 1 0 19872 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_208
timestamp 1644511149
transform 1 0 20240 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_211
timestamp 1644511149
transform 1 0 20516 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 1644511149
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_225
timestamp 1644511149
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_237
timestamp 1644511149
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_249
timestamp 1644511149
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_261
timestamp 1644511149
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_273
timestamp 1644511149
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1644511149
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_281
timestamp 1644511149
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_293
timestamp 1644511149
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_305
timestamp 1644511149
transform 1 0 29164 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_317
timestamp 1644511149
transform 1 0 30268 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_329
timestamp 1644511149
transform 1 0 31372 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_335
timestamp 1644511149
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_337
timestamp 1644511149
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_349
timestamp 1644511149
transform 1 0 33212 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_357
timestamp 1644511149
transform 1 0 33948 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_362
timestamp 1644511149
transform 1 0 34408 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_42_3
timestamp 1644511149
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_15
timestamp 1644511149
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1644511149
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_29
timestamp 1644511149
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_41
timestamp 1644511149
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_53
timestamp 1644511149
transform 1 0 5980 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_57
timestamp 1644511149
transform 1 0 6348 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_69
timestamp 1644511149
transform 1 0 7452 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_81
timestamp 1644511149
transform 1 0 8556 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_85
timestamp 1644511149
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_97
timestamp 1644511149
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_109
timestamp 1644511149
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_121
timestamp 1644511149
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_133
timestamp 1644511149
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1644511149
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_141
timestamp 1644511149
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_153
timestamp 1644511149
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_165
timestamp 1644511149
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_177
timestamp 1644511149
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_189
timestamp 1644511149
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1644511149
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_200
timestamp 1644511149
transform 1 0 19504 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_209
timestamp 1644511149
transform 1 0 20332 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_214
timestamp 1644511149
transform 1 0 20792 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_42_218
timestamp 1644511149
transform 1 0 21160 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_230
timestamp 1644511149
transform 1 0 22264 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_242
timestamp 1644511149
transform 1 0 23368 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_250
timestamp 1644511149
transform 1 0 24104 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_42_253
timestamp 1644511149
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_265
timestamp 1644511149
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_277
timestamp 1644511149
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_289
timestamp 1644511149
transform 1 0 27692 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_301
timestamp 1644511149
transform 1 0 28796 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 1644511149
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_309
timestamp 1644511149
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_321
timestamp 1644511149
transform 1 0 30636 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_333
timestamp 1644511149
transform 1 0 31740 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_345
timestamp 1644511149
transform 1 0 32844 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_357
timestamp 1644511149
transform 1 0 33948 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_362
timestamp 1644511149
transform 1 0 34408 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_43_3
timestamp 1644511149
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_15
timestamp 1644511149
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_27
timestamp 1644511149
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_39
timestamp 1644511149
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1644511149
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1644511149
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_57
timestamp 1644511149
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_69
timestamp 1644511149
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_81
timestamp 1644511149
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_93
timestamp 1644511149
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1644511149
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1644511149
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_113
timestamp 1644511149
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_125
timestamp 1644511149
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_137
timestamp 1644511149
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_149
timestamp 1644511149
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_161
timestamp 1644511149
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1644511149
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_169
timestamp 1644511149
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_185
timestamp 1644511149
transform 1 0 18124 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_191
timestamp 1644511149
transform 1 0 18676 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_195
timestamp 1644511149
transform 1 0 19044 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_202
timestamp 1644511149
transform 1 0 19688 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_212
timestamp 1644511149
transform 1 0 20608 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_220
timestamp 1644511149
transform 1 0 21344 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_227
timestamp 1644511149
transform 1 0 21988 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_239
timestamp 1644511149
transform 1 0 23092 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_251
timestamp 1644511149
transform 1 0 24196 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_263
timestamp 1644511149
transform 1 0 25300 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_275
timestamp 1644511149
transform 1 0 26404 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1644511149
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_281
timestamp 1644511149
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_293
timestamp 1644511149
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_305
timestamp 1644511149
transform 1 0 29164 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_317
timestamp 1644511149
transform 1 0 30268 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_329
timestamp 1644511149
transform 1 0 31372 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1644511149
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_337
timestamp 1644511149
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_349
timestamp 1644511149
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_43_361
timestamp 1644511149
transform 1 0 34316 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_44_6
timestamp 1644511149
transform 1 0 1656 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_44_10
timestamp 1644511149
transform 1 0 2024 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_22
timestamp 1644511149
transform 1 0 3128 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_44_29
timestamp 1644511149
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_41
timestamp 1644511149
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_53
timestamp 1644511149
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_65
timestamp 1644511149
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1644511149
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1644511149
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_85
timestamp 1644511149
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_97
timestamp 1644511149
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_109
timestamp 1644511149
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_121
timestamp 1644511149
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 1644511149
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1644511149
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_141
timestamp 1644511149
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_153
timestamp 1644511149
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_165
timestamp 1644511149
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_177
timestamp 1644511149
transform 1 0 17388 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_44_187
timestamp 1644511149
transform 1 0 18308 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_194
timestamp 1644511149
transform 1 0 18952 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_44_197
timestamp 1644511149
transform 1 0 19228 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_44_209
timestamp 1644511149
transform 1 0 20332 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_217
timestamp 1644511149
transform 1 0 21068 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_224
timestamp 1644511149
transform 1 0 21712 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_44_228
timestamp 1644511149
transform 1 0 22080 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_240
timestamp 1644511149
transform 1 0 23184 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_253
timestamp 1644511149
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_265
timestamp 1644511149
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_277
timestamp 1644511149
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_289
timestamp 1644511149
transform 1 0 27692 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_301
timestamp 1644511149
transform 1 0 28796 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 1644511149
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_309
timestamp 1644511149
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_321
timestamp 1644511149
transform 1 0 30636 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_333
timestamp 1644511149
transform 1 0 31740 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_345
timestamp 1644511149
transform 1 0 32844 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_353
timestamp 1644511149
transform 1 0 33580 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_357
timestamp 1644511149
transform 1 0 33948 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_362
timestamp 1644511149
transform 1 0 34408 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_45_3
timestamp 1644511149
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_15
timestamp 1644511149
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_27
timestamp 1644511149
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_39
timestamp 1644511149
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1644511149
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1644511149
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_57
timestamp 1644511149
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_69
timestamp 1644511149
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_81
timestamp 1644511149
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_93
timestamp 1644511149
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 1644511149
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1644511149
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_113
timestamp 1644511149
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_125
timestamp 1644511149
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_137
timestamp 1644511149
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_149
timestamp 1644511149
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_161
timestamp 1644511149
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1644511149
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_169
timestamp 1644511149
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_185
timestamp 1644511149
transform 1 0 18124 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_189
timestamp 1644511149
transform 1 0 18492 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_192
timestamp 1644511149
transform 1 0 18768 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_45_196
timestamp 1644511149
transform 1 0 19136 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_45_207
timestamp 1644511149
transform 1 0 20148 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_216
timestamp 1644511149
transform 1 0 20976 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_45_221
timestamp 1644511149
transform 1 0 21436 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_45_227
timestamp 1644511149
transform 1 0 21988 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_45_231
timestamp 1644511149
transform 1 0 22356 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_243
timestamp 1644511149
transform 1 0 23460 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_255
timestamp 1644511149
transform 1 0 24564 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_267
timestamp 1644511149
transform 1 0 25668 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 1644511149
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_281
timestamp 1644511149
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_293
timestamp 1644511149
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_305
timestamp 1644511149
transform 1 0 29164 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_317
timestamp 1644511149
transform 1 0 30268 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_329
timestamp 1644511149
transform 1 0 31372 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 1644511149
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_337
timestamp 1644511149
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_349
timestamp 1644511149
transform 1 0 33212 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_353
timestamp 1644511149
transform 1 0 33580 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_356
timestamp 1644511149
transform 1 0 33856 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_362
timestamp 1644511149
transform 1 0 34408 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_46_3
timestamp 1644511149
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_15
timestamp 1644511149
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1644511149
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_29
timestamp 1644511149
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_41
timestamp 1644511149
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_53
timestamp 1644511149
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_65
timestamp 1644511149
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1644511149
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1644511149
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_85
timestamp 1644511149
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_97
timestamp 1644511149
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_109
timestamp 1644511149
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_121
timestamp 1644511149
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 1644511149
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1644511149
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_141
timestamp 1644511149
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_153
timestamp 1644511149
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_165
timestamp 1644511149
transform 1 0 16284 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_177
timestamp 1644511149
transform 1 0 17388 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_189
timestamp 1644511149
transform 1 0 18492 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1644511149
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_199
timestamp 1644511149
transform 1 0 19412 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_208
timestamp 1644511149
transform 1 0 20240 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_213
timestamp 1644511149
transform 1 0 20700 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_217
timestamp 1644511149
transform 1 0 21068 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_221
timestamp 1644511149
transform 1 0 21436 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_46_225
timestamp 1644511149
transform 1 0 21804 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_237
timestamp 1644511149
transform 1 0 22908 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_249
timestamp 1644511149
transform 1 0 24012 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_253
timestamp 1644511149
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_265
timestamp 1644511149
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_277
timestamp 1644511149
transform 1 0 26588 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_289
timestamp 1644511149
transform 1 0 27692 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_301
timestamp 1644511149
transform 1 0 28796 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_307
timestamp 1644511149
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_309
timestamp 1644511149
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_321
timestamp 1644511149
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_333
timestamp 1644511149
transform 1 0 31740 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_345
timestamp 1644511149
transform 1 0 32844 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_357
timestamp 1644511149
transform 1 0 33948 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1644511149
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_7
timestamp 1644511149
transform 1 0 1748 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_47_11
timestamp 1644511149
transform 1 0 2116 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_23
timestamp 1644511149
transform 1 0 3220 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_35
timestamp 1644511149
transform 1 0 4324 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_47
timestamp 1644511149
transform 1 0 5428 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1644511149
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_57
timestamp 1644511149
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_69
timestamp 1644511149
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_81
timestamp 1644511149
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_93
timestamp 1644511149
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_105
timestamp 1644511149
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1644511149
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_113
timestamp 1644511149
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_125
timestamp 1644511149
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_137
timestamp 1644511149
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_149
timestamp 1644511149
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_161
timestamp 1644511149
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1644511149
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_169
timestamp 1644511149
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_181
timestamp 1644511149
transform 1 0 17756 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_193
timestamp 1644511149
transform 1 0 18860 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_47_205
timestamp 1644511149
transform 1 0 19964 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_47_210
timestamp 1644511149
transform 1 0 20424 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_222
timestamp 1644511149
transform 1 0 21528 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_47_225
timestamp 1644511149
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_237
timestamp 1644511149
transform 1 0 22908 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_249
timestamp 1644511149
transform 1 0 24012 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_261
timestamp 1644511149
transform 1 0 25116 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_273
timestamp 1644511149
transform 1 0 26220 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_279
timestamp 1644511149
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_281
timestamp 1644511149
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_293
timestamp 1644511149
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_305
timestamp 1644511149
transform 1 0 29164 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_317
timestamp 1644511149
transform 1 0 30268 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_323
timestamp 1644511149
transform 1 0 30820 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_327
timestamp 1644511149
transform 1 0 31188 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_335
timestamp 1644511149
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_337
timestamp 1644511149
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_349
timestamp 1644511149
transform 1 0 33212 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_357
timestamp 1644511149
transform 1 0 33948 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_362
timestamp 1644511149
transform 1 0 34408 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_48_3
timestamp 1644511149
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_15
timestamp 1644511149
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1644511149
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_29
timestamp 1644511149
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_41
timestamp 1644511149
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_53
timestamp 1644511149
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_65
timestamp 1644511149
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1644511149
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1644511149
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_85
timestamp 1644511149
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_97
timestamp 1644511149
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_109
timestamp 1644511149
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_121
timestamp 1644511149
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_133
timestamp 1644511149
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1644511149
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_141
timestamp 1644511149
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_153
timestamp 1644511149
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_165
timestamp 1644511149
transform 1 0 16284 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_177
timestamp 1644511149
transform 1 0 17388 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_189
timestamp 1644511149
transform 1 0 18492 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1644511149
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_197
timestamp 1644511149
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_209
timestamp 1644511149
transform 1 0 20332 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_221
timestamp 1644511149
transform 1 0 21436 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_233
timestamp 1644511149
transform 1 0 22540 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_245
timestamp 1644511149
transform 1 0 23644 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1644511149
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_253
timestamp 1644511149
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_265
timestamp 1644511149
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_277
timestamp 1644511149
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_289
timestamp 1644511149
transform 1 0 27692 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_301
timestamp 1644511149
transform 1 0 28796 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_307
timestamp 1644511149
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_309
timestamp 1644511149
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_321
timestamp 1644511149
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_333
timestamp 1644511149
transform 1 0 31740 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_345
timestamp 1644511149
transform 1 0 32844 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_353
timestamp 1644511149
transform 1 0 33580 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_48_358
timestamp 1644511149
transform 1 0 34040 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_49_3
timestamp 1644511149
transform 1 0 1380 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_9
timestamp 1644511149
transform 1 0 1932 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_49_13
timestamp 1644511149
transform 1 0 2300 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_25
timestamp 1644511149
transform 1 0 3404 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_37
timestamp 1644511149
transform 1 0 4508 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_49
timestamp 1644511149
transform 1 0 5612 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1644511149
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_57
timestamp 1644511149
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_69
timestamp 1644511149
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_81
timestamp 1644511149
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_93
timestamp 1644511149
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 1644511149
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1644511149
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_113
timestamp 1644511149
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_125
timestamp 1644511149
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_137
timestamp 1644511149
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_149
timestamp 1644511149
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_161
timestamp 1644511149
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1644511149
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_169
timestamp 1644511149
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_181
timestamp 1644511149
transform 1 0 17756 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_193
timestamp 1644511149
transform 1 0 18860 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_205
timestamp 1644511149
transform 1 0 19964 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_217
timestamp 1644511149
transform 1 0 21068 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 1644511149
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_225
timestamp 1644511149
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_237
timestamp 1644511149
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_249
timestamp 1644511149
transform 1 0 24012 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_261
timestamp 1644511149
transform 1 0 25116 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_273
timestamp 1644511149
transform 1 0 26220 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 1644511149
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_281
timestamp 1644511149
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_293
timestamp 1644511149
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_305
timestamp 1644511149
transform 1 0 29164 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_317
timestamp 1644511149
transform 1 0 30268 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_329
timestamp 1644511149
transform 1 0 31372 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 1644511149
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_337
timestamp 1644511149
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_349
timestamp 1644511149
transform 1 0 33212 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_356
timestamp 1644511149
transform 1 0 33856 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_362
timestamp 1644511149
transform 1 0 34408 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_7
timestamp 1644511149
transform 1 0 1748 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_11
timestamp 1644511149
transform 1 0 2116 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_50_15
timestamp 1644511149
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1644511149
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_29
timestamp 1644511149
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_41
timestamp 1644511149
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_53
timestamp 1644511149
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_65
timestamp 1644511149
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1644511149
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1644511149
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_85
timestamp 1644511149
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_97
timestamp 1644511149
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_109
timestamp 1644511149
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_121
timestamp 1644511149
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 1644511149
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1644511149
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_141
timestamp 1644511149
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_153
timestamp 1644511149
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_165
timestamp 1644511149
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_177
timestamp 1644511149
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_189
timestamp 1644511149
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1644511149
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_197
timestamp 1644511149
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_209
timestamp 1644511149
transform 1 0 20332 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_221
timestamp 1644511149
transform 1 0 21436 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_233
timestamp 1644511149
transform 1 0 22540 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_245
timestamp 1644511149
transform 1 0 23644 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 1644511149
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_253
timestamp 1644511149
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_265
timestamp 1644511149
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_277
timestamp 1644511149
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_289
timestamp 1644511149
transform 1 0 27692 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_301
timestamp 1644511149
transform 1 0 28796 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_307
timestamp 1644511149
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_309
timestamp 1644511149
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_321
timestamp 1644511149
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_333
timestamp 1644511149
transform 1 0 31740 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_345
timestamp 1644511149
transform 1 0 32844 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_353
timestamp 1644511149
transform 1 0 33580 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_357
timestamp 1644511149
transform 1 0 33948 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_362
timestamp 1644511149
transform 1 0 34408 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_51_13
timestamp 1644511149
transform 1 0 2300 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_25
timestamp 1644511149
transform 1 0 3404 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_37
timestamp 1644511149
transform 1 0 4508 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_49
timestamp 1644511149
transform 1 0 5612 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1644511149
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_57
timestamp 1644511149
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_69
timestamp 1644511149
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_81
timestamp 1644511149
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_93
timestamp 1644511149
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1644511149
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1644511149
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_113
timestamp 1644511149
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_125
timestamp 1644511149
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_137
timestamp 1644511149
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_149
timestamp 1644511149
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_161
timestamp 1644511149
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1644511149
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_169
timestamp 1644511149
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_181
timestamp 1644511149
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_193
timestamp 1644511149
transform 1 0 18860 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_205
timestamp 1644511149
transform 1 0 19964 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_217
timestamp 1644511149
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1644511149
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_225
timestamp 1644511149
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_237
timestamp 1644511149
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_249
timestamp 1644511149
transform 1 0 24012 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_261
timestamp 1644511149
transform 1 0 25116 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_273
timestamp 1644511149
transform 1 0 26220 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1644511149
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_281
timestamp 1644511149
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_293
timestamp 1644511149
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_305
timestamp 1644511149
transform 1 0 29164 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_317
timestamp 1644511149
transform 1 0 30268 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_329
timestamp 1644511149
transform 1 0 31372 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_335
timestamp 1644511149
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_337
timestamp 1644511149
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_349
timestamp 1644511149
transform 1 0 33212 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_353
timestamp 1644511149
transform 1 0 33580 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_357
timestamp 1644511149
transform 1 0 33948 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_362
timestamp 1644511149
transform 1 0 34408 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_7
timestamp 1644511149
transform 1 0 1748 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_52_11
timestamp 1644511149
transform 1 0 2116 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_23
timestamp 1644511149
transform 1 0 3220 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1644511149
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_29
timestamp 1644511149
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_41
timestamp 1644511149
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_53
timestamp 1644511149
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_65
timestamp 1644511149
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1644511149
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1644511149
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_85
timestamp 1644511149
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_97
timestamp 1644511149
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_109
timestamp 1644511149
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_121
timestamp 1644511149
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1644511149
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1644511149
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_141
timestamp 1644511149
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_153
timestamp 1644511149
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_165
timestamp 1644511149
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_177
timestamp 1644511149
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_189
timestamp 1644511149
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1644511149
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_197
timestamp 1644511149
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_209
timestamp 1644511149
transform 1 0 20332 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_221
timestamp 1644511149
transform 1 0 21436 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_233
timestamp 1644511149
transform 1 0 22540 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_245
timestamp 1644511149
transform 1 0 23644 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1644511149
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_253
timestamp 1644511149
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_265
timestamp 1644511149
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_277
timestamp 1644511149
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_289
timestamp 1644511149
transform 1 0 27692 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_301
timestamp 1644511149
transform 1 0 28796 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1644511149
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_309
timestamp 1644511149
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_321
timestamp 1644511149
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_333
timestamp 1644511149
transform 1 0 31740 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_345
timestamp 1644511149
transform 1 0 32844 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_351
timestamp 1644511149
transform 1 0 33396 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_362
timestamp 1644511149
transform 1 0 34408 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_53_5
timestamp 1644511149
transform 1 0 1564 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_17
timestamp 1644511149
transform 1 0 2668 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_29
timestamp 1644511149
transform 1 0 3772 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_41
timestamp 1644511149
transform 1 0 4876 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_53_53
timestamp 1644511149
transform 1 0 5980 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_53_57
timestamp 1644511149
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_69
timestamp 1644511149
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_81
timestamp 1644511149
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_93
timestamp 1644511149
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1644511149
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1644511149
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_113
timestamp 1644511149
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_125
timestamp 1644511149
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_137
timestamp 1644511149
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_149
timestamp 1644511149
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_161
timestamp 1644511149
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1644511149
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_169
timestamp 1644511149
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_185
timestamp 1644511149
transform 1 0 18124 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_197
timestamp 1644511149
transform 1 0 19228 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_209
timestamp 1644511149
transform 1 0 20332 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_53_221
timestamp 1644511149
transform 1 0 21436 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_53_225
timestamp 1644511149
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_237
timestamp 1644511149
transform 1 0 22908 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_249
timestamp 1644511149
transform 1 0 24012 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_261
timestamp 1644511149
transform 1 0 25116 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_273
timestamp 1644511149
transform 1 0 26220 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1644511149
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_281
timestamp 1644511149
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_293
timestamp 1644511149
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_305
timestamp 1644511149
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_317
timestamp 1644511149
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_329
timestamp 1644511149
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1644511149
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_337
timestamp 1644511149
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_349
timestamp 1644511149
transform 1 0 33212 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_353
timestamp 1644511149
transform 1 0 33580 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_357
timestamp 1644511149
transform 1 0 33948 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_362
timestamp 1644511149
transform 1 0 34408 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_7
timestamp 1644511149
transform 1 0 1748 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_13
timestamp 1644511149
transform 1 0 2300 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_17
timestamp 1644511149
transform 1 0 2668 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_54_21
timestamp 1644511149
transform 1 0 3036 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1644511149
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_29
timestamp 1644511149
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_41
timestamp 1644511149
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_53
timestamp 1644511149
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_65
timestamp 1644511149
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1644511149
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1644511149
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_85
timestamp 1644511149
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_97
timestamp 1644511149
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_109
timestamp 1644511149
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_121
timestamp 1644511149
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1644511149
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1644511149
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_141
timestamp 1644511149
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_153
timestamp 1644511149
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_165
timestamp 1644511149
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_177
timestamp 1644511149
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_189
timestamp 1644511149
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 1644511149
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_197
timestamp 1644511149
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_209
timestamp 1644511149
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_221
timestamp 1644511149
transform 1 0 21436 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_233
timestamp 1644511149
transform 1 0 22540 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_245
timestamp 1644511149
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1644511149
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_253
timestamp 1644511149
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_265
timestamp 1644511149
transform 1 0 25484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_277
timestamp 1644511149
transform 1 0 26588 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_289
timestamp 1644511149
transform 1 0 27692 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_301
timestamp 1644511149
transform 1 0 28796 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1644511149
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_309
timestamp 1644511149
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_321
timestamp 1644511149
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_333
timestamp 1644511149
transform 1 0 31740 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_343
timestamp 1644511149
transform 1 0 32660 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_347
timestamp 1644511149
transform 1 0 33028 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_351
timestamp 1644511149
transform 1 0 33396 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_356
timestamp 1644511149
transform 1 0 33856 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_362
timestamp 1644511149
transform 1 0 34408 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_13
timestamp 1644511149
transform 1 0 2300 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_19
timestamp 1644511149
transform 1 0 2852 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_55_23
timestamp 1644511149
transform 1 0 3220 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_35
timestamp 1644511149
transform 1 0 4324 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_47
timestamp 1644511149
transform 1 0 5428 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1644511149
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_57
timestamp 1644511149
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_69
timestamp 1644511149
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_81
timestamp 1644511149
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_93
timestamp 1644511149
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1644511149
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1644511149
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_113
timestamp 1644511149
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_125
timestamp 1644511149
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_137
timestamp 1644511149
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_149
timestamp 1644511149
transform 1 0 14812 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_55_158
timestamp 1644511149
transform 1 0 15640 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_166
timestamp 1644511149
transform 1 0 16376 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_55_169
timestamp 1644511149
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_181
timestamp 1644511149
transform 1 0 17756 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_186
timestamp 1644511149
transform 1 0 18216 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_192
timestamp 1644511149
transform 1 0 18768 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_55_196
timestamp 1644511149
transform 1 0 19136 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_208
timestamp 1644511149
transform 1 0 20240 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_220
timestamp 1644511149
transform 1 0 21344 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_225
timestamp 1644511149
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_237
timestamp 1644511149
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_249
timestamp 1644511149
transform 1 0 24012 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_261
timestamp 1644511149
transform 1 0 25116 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_273
timestamp 1644511149
transform 1 0 26220 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 1644511149
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_281
timestamp 1644511149
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_293
timestamp 1644511149
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_305
timestamp 1644511149
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_317
timestamp 1644511149
transform 1 0 30268 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_55_329
timestamp 1644511149
transform 1 0 31372 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_55_334
timestamp 1644511149
transform 1 0 31832 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_337
timestamp 1644511149
transform 1 0 32108 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_341
timestamp 1644511149
transform 1 0 32476 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_345
timestamp 1644511149
transform 1 0 32844 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_350
timestamp 1644511149
transform 1 0 33304 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_356
timestamp 1644511149
transform 1 0 33856 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_362
timestamp 1644511149
transform 1 0 34408 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_3
timestamp 1644511149
transform 1 0 1380 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_9
timestamp 1644511149
transform 1 0 1932 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_15
timestamp 1644511149
transform 1 0 2484 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_19
timestamp 1644511149
transform 1 0 2852 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_56_25
timestamp 1644511149
transform 1 0 3404 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_56_29
timestamp 1644511149
transform 1 0 3772 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_35
timestamp 1644511149
transform 1 0 4324 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_38
timestamp 1644511149
transform 1 0 4600 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_46
timestamp 1644511149
transform 1 0 5336 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_50
timestamp 1644511149
transform 1 0 5704 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_56
timestamp 1644511149
transform 1 0 6256 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_56_60
timestamp 1644511149
transform 1 0 6624 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_72
timestamp 1644511149
transform 1 0 7728 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_82
timestamp 1644511149
transform 1 0 8648 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_85
timestamp 1644511149
transform 1 0 8924 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_90
timestamp 1644511149
transform 1 0 9384 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_56_94
timestamp 1644511149
transform 1 0 9752 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_102
timestamp 1644511149
transform 1 0 10488 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_106
timestamp 1644511149
transform 1 0 10856 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_111
timestamp 1644511149
transform 1 0 11316 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_56_115
timestamp 1644511149
transform 1 0 11684 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_127
timestamp 1644511149
transform 1 0 12788 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1644511149
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_141
timestamp 1644511149
transform 1 0 14076 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_145
timestamp 1644511149
transform 1 0 14444 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_148
timestamp 1644511149
transform 1 0 14720 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_160
timestamp 1644511149
transform 1 0 15824 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_168
timestamp 1644511149
transform 1 0 16560 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_173
timestamp 1644511149
transform 1 0 17020 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_180
timestamp 1644511149
transform 1 0 17664 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_186
timestamp 1644511149
transform 1 0 18216 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_192
timestamp 1644511149
transform 1 0 18768 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_201
timestamp 1644511149
transform 1 0 19596 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_213
timestamp 1644511149
transform 1 0 20700 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_221
timestamp 1644511149
transform 1 0 21436 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_224
timestamp 1644511149
transform 1 0 21712 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_56_229
timestamp 1644511149
transform 1 0 22172 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_241
timestamp 1644511149
transform 1 0 23276 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_56_249
timestamp 1644511149
transform 1 0 24012 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_56_253
timestamp 1644511149
transform 1 0 24380 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_56_259
timestamp 1644511149
transform 1 0 24932 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_56_266
timestamp 1644511149
transform 1 0 25576 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_278
timestamp 1644511149
transform 1 0 26680 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_282
timestamp 1644511149
transform 1 0 27048 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_287
timestamp 1644511149
transform 1 0 27508 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_56_292
timestamp 1644511149
transform 1 0 27968 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_56_302
timestamp 1644511149
transform 1 0 28888 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_56_309
timestamp 1644511149
transform 1 0 29532 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_315
timestamp 1644511149
transform 1 0 30084 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_56_318
timestamp 1644511149
transform 1 0 30360 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_56_323
timestamp 1644511149
transform 1 0 30820 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_335
timestamp 1644511149
transform 1 0 31924 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_56_343
timestamp 1644511149
transform 1 0 32660 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_56_350
timestamp 1644511149
transform 1 0 33304 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_356
timestamp 1644511149
transform 1 0 33856 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_362
timestamp 1644511149
transform 1 0 34408 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_13
timestamp 1644511149
transform 1 0 2300 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_21
timestamp 1644511149
transform 1 0 3036 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_57_25
timestamp 1644511149
transform 1 0 3404 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_57_29
timestamp 1644511149
transform 1 0 3772 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_57_35
timestamp 1644511149
transform 1 0 4324 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_57_48
timestamp 1644511149
transform 1 0 5520 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_54
timestamp 1644511149
transform 1 0 6072 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_57
timestamp 1644511149
transform 1 0 6348 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_57_63
timestamp 1644511149
transform 1 0 6900 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_71
timestamp 1644511149
transform 1 0 7636 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_77
timestamp 1644511149
transform 1 0 8188 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_57_81
timestamp 1644511149
transform 1 0 8556 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_57_85
timestamp 1644511149
transform 1 0 8924 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_57_91
timestamp 1644511149
transform 1 0 9476 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_57_98
timestamp 1644511149
transform 1 0 10120 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_110
timestamp 1644511149
transform 1 0 11224 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_113
timestamp 1644511149
transform 1 0 11500 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_118
timestamp 1644511149
transform 1 0 11960 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_57_122
timestamp 1644511149
transform 1 0 12328 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_134
timestamp 1644511149
transform 1 0 13432 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_138
timestamp 1644511149
transform 1 0 13800 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_145
timestamp 1644511149
transform 1 0 14444 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_150
timestamp 1644511149
transform 1 0 14904 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_154
timestamp 1644511149
transform 1 0 15272 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_166
timestamp 1644511149
transform 1 0 16376 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_169
timestamp 1644511149
transform 1 0 16652 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_175
timestamp 1644511149
transform 1 0 17204 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_57_179
timestamp 1644511149
transform 1 0 17572 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_57_189
timestamp 1644511149
transform 1 0 18492 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_57_194
timestamp 1644511149
transform 1 0 18952 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_197
timestamp 1644511149
transform 1 0 19228 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_57_209
timestamp 1644511149
transform 1 0 20332 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_57_222
timestamp 1644511149
transform 1 0 21528 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_228
timestamp 1644511149
transform 1 0 22080 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_232
timestamp 1644511149
transform 1 0 22448 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_236
timestamp 1644511149
transform 1 0 22816 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_239
timestamp 1644511149
transform 1 0 23092 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_244
timestamp 1644511149
transform 1 0 23552 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_250
timestamp 1644511149
transform 1 0 24104 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_263
timestamp 1644511149
transform 1 0 25300 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_267
timestamp 1644511149
transform 1 0 25668 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_57_273
timestamp 1644511149
transform 1 0 26220 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_57_278
timestamp 1644511149
transform 1 0 26680 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_291
timestamp 1644511149
transform 1 0 27876 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_295
timestamp 1644511149
transform 1 0 28244 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_300
timestamp 1644511149
transform 1 0 28704 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_306
timestamp 1644511149
transform 1 0 29256 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_309
timestamp 1644511149
transform 1 0 29532 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_57_315
timestamp 1644511149
transform 1 0 30084 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_57_328
timestamp 1644511149
transform 1 0 31280 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_334
timestamp 1644511149
transform 1 0 31832 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_337
timestamp 1644511149
transform 1 0 32108 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_57_343
timestamp 1644511149
transform 1 0 32660 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_57_350
timestamp 1644511149
transform 1 0 33304 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_362
timestamp 1644511149
transform 1 0 34408 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1644511149
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1644511149
transform -1 0 34868 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1644511149
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1644511149
transform -1 0 34868 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1644511149
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1644511149
transform -1 0 34868 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1644511149
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1644511149
transform -1 0 34868 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1644511149
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1644511149
transform -1 0 34868 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1644511149
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1644511149
transform -1 0 34868 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1644511149
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1644511149
transform -1 0 34868 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1644511149
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1644511149
transform -1 0 34868 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1644511149
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1644511149
transform -1 0 34868 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1644511149
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1644511149
transform -1 0 34868 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1644511149
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1644511149
transform -1 0 34868 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1644511149
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1644511149
transform -1 0 34868 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1644511149
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1644511149
transform -1 0 34868 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1644511149
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1644511149
transform -1 0 34868 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1644511149
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1644511149
transform -1 0 34868 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1644511149
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1644511149
transform -1 0 34868 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1644511149
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1644511149
transform -1 0 34868 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1644511149
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1644511149
transform -1 0 34868 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1644511149
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1644511149
transform -1 0 34868 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1644511149
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1644511149
transform -1 0 34868 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1644511149
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1644511149
transform -1 0 34868 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1644511149
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1644511149
transform -1 0 34868 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1644511149
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1644511149
transform -1 0 34868 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1644511149
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1644511149
transform -1 0 34868 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1644511149
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1644511149
transform -1 0 34868 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1644511149
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1644511149
transform -1 0 34868 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1644511149
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1644511149
transform -1 0 34868 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1644511149
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1644511149
transform -1 0 34868 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1644511149
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1644511149
transform -1 0 34868 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1644511149
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1644511149
transform -1 0 34868 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1644511149
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1644511149
transform -1 0 34868 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1644511149
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1644511149
transform -1 0 34868 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1644511149
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1644511149
transform -1 0 34868 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1644511149
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1644511149
transform -1 0 34868 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1644511149
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1644511149
transform -1 0 34868 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1644511149
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1644511149
transform -1 0 34868 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1644511149
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1644511149
transform -1 0 34868 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1644511149
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1644511149
transform -1 0 34868 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1644511149
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1644511149
transform -1 0 34868 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1644511149
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1644511149
transform -1 0 34868 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1644511149
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1644511149
transform -1 0 34868 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1644511149
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1644511149
transform -1 0 34868 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1644511149
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1644511149
transform -1 0 34868 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1644511149
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1644511149
transform -1 0 34868 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1644511149
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1644511149
transform -1 0 34868 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1644511149
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1644511149
transform -1 0 34868 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1644511149
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1644511149
transform -1 0 34868 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1644511149
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1644511149
transform -1 0 34868 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1644511149
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1644511149
transform -1 0 34868 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1644511149
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1644511149
transform -1 0 34868 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1644511149
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1644511149
transform -1 0 34868 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1644511149
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1644511149
transform -1 0 34868 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1644511149
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1644511149
transform -1 0 34868 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1644511149
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1644511149
transform -1 0 34868 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1644511149
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1644511149
transform -1 0 34868 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1644511149
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1644511149
transform -1 0 34868 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1644511149
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1644511149
transform -1 0 34868 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1644511149
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1644511149
transform -1 0 34868 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1644511149
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1644511149
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1644511149
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1644511149
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1644511149
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1644511149
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1644511149
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1644511149
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1644511149
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1644511149
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1644511149
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1644511149
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1644511149
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1644511149
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1644511149
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1644511149
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1644511149
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1644511149
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1644511149
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1644511149
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1644511149
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1644511149
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1644511149
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1644511149
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1644511149
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1644511149
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1644511149
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1644511149
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1644511149
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1644511149
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1644511149
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1644511149
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1644511149
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1644511149
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1644511149
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1644511149
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1644511149
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1644511149
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1644511149
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1644511149
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1644511149
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1644511149
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1644511149
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1644511149
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1644511149
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1644511149
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1644511149
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1644511149
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1644511149
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1644511149
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1644511149
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1644511149
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1644511149
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1644511149
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1644511149
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1644511149
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1644511149
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1644511149
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1644511149
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1644511149
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1644511149
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1644511149
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1644511149
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1644511149
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1644511149
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1644511149
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1644511149
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1644511149
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1644511149
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1644511149
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1644511149
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1644511149
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1644511149
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1644511149
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1644511149
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1644511149
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1644511149
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1644511149
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1644511149
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1644511149
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1644511149
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1644511149
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1644511149
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1644511149
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1644511149
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1644511149
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1644511149
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1644511149
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1644511149
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1644511149
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1644511149
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1644511149
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1644511149
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1644511149
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1644511149
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1644511149
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1644511149
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1644511149
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1644511149
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1644511149
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1644511149
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1644511149
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1644511149
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1644511149
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1644511149
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1644511149
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1644511149
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1644511149
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1644511149
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1644511149
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1644511149
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1644511149
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1644511149
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1644511149
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1644511149
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1644511149
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1644511149
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1644511149
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1644511149
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1644511149
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1644511149
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1644511149
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1644511149
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1644511149
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1644511149
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1644511149
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1644511149
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1644511149
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1644511149
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1644511149
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1644511149
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1644511149
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1644511149
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1644511149
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1644511149
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1644511149
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1644511149
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1644511149
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1644511149
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1644511149
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1644511149
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1644511149
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1644511149
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1644511149
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1644511149
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1644511149
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1644511149
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1644511149
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1644511149
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1644511149
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1644511149
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1644511149
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1644511149
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1644511149
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1644511149
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1644511149
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1644511149
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1644511149
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1644511149
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1644511149
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1644511149
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1644511149
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1644511149
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1644511149
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1644511149
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1644511149
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1644511149
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1644511149
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1644511149
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1644511149
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1644511149
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1644511149
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1644511149
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1644511149
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1644511149
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1644511149
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1644511149
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1644511149
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1644511149
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1644511149
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1644511149
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1644511149
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1644511149
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1644511149
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1644511149
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1644511149
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1644511149
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1644511149
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1644511149
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1644511149
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1644511149
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1644511149
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1644511149
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1644511149
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1644511149
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1644511149
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1644511149
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1644511149
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1644511149
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1644511149
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1644511149
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1644511149
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1644511149
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1644511149
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1644511149
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1644511149
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1644511149
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1644511149
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1644511149
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1644511149
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1644511149
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1644511149
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1644511149
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1644511149
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1644511149
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1644511149
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1644511149
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1644511149
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1644511149
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1644511149
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1644511149
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1644511149
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1644511149
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1644511149
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1644511149
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1644511149
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1644511149
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1644511149
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1644511149
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1644511149
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1644511149
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1644511149
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1644511149
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1644511149
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1644511149
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1644511149
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1644511149
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1644511149
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1644511149
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1644511149
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1644511149
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1644511149
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1644511149
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1644511149
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1644511149
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1644511149
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1644511149
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1644511149
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1644511149
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1644511149
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1644511149
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1644511149
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1644511149
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1644511149
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1644511149
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1644511149
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1644511149
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1644511149
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1644511149
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1644511149
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1644511149
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1644511149
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1644511149
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1644511149
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1644511149
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1644511149
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1644511149
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1644511149
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1644511149
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1644511149
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1644511149
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1644511149
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1644511149
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1644511149
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1644511149
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1644511149
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1644511149
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1644511149
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1644511149
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1644511149
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1644511149
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1644511149
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1644511149
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1644511149
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1644511149
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1644511149
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1644511149
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1644511149
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1644511149
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1644511149
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1644511149
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1644511149
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1644511149
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1644511149
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1644511149
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1644511149
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1644511149
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1644511149
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1644511149
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1644511149
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1644511149
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1644511149
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1644511149
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1644511149
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1644511149
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1644511149
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1644511149
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1644511149
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1644511149
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1644511149
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1644511149
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1644511149
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1644511149
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1644511149
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1644511149
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1644511149
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1644511149
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1644511149
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1644511149
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1644511149
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1644511149
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1644511149
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1644511149
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1644511149
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1644511149
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1644511149
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1644511149
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1644511149
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1644511149
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1644511149
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1644511149
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1644511149
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1644511149
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1644511149
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1644511149
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1644511149
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1644511149
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1644511149
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1644511149
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1644511149
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1644511149
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1644511149
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1644511149
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1644511149
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1644511149
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1644511149
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1644511149
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1644511149
transform 1 0 3680 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1644511149
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1644511149
transform 1 0 8832 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1644511149
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1644511149
transform 1 0 13984 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1644511149
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1644511149
transform 1 0 19136 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1644511149
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1644511149
transform 1 0 24288 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1644511149
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1644511149
transform 1 0 29440 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1644511149
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _011_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 18676 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _012_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 20976 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _013_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20516 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _014_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 20700 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _015_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20516 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a311o_2  _016_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19504 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__or2b_1  _017_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 21344 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _018_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 21712 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _019_
timestamp 1644511149
transform -1 0 21436 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _020_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19596 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _021_
timestamp 1644511149
transform -1 0 20332 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_2  _022_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 20608 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _023_
timestamp 1644511149
transform 1 0 19228 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_2  _024_
timestamp 1644511149
transform 1 0 19412 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _025_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 29624 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _026_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 29532 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _027_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17756 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _028_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 8924 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _029_
timestamp 1644511149
transform -1 0 18676 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _030_
timestamp 1644511149
transform 1 0 17848 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _031_
timestamp 1644511149
transform -1 0 18216 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _032_
timestamp 1644511149
transform 1 0 17848 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _033_
timestamp 1644511149
transform -1 0 33856 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _034_
timestamp 1644511149
transform -1 0 17664 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _035_
timestamp 1644511149
transform 1 0 17204 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _036_
timestamp 1644511149
transform -1 0 18216 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _037_
timestamp 1644511149
transform 1 0 17848 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _038_
timestamp 1644511149
transform -1 0 18216 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _039_
timestamp 1644511149
transform 1 0 18860 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _040_
timestamp 1644511149
transform -1 0 18768 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _041_
timestamp 1644511149
transform 1 0 7084 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _042_
timestamp 1644511149
transform -1 0 18124 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _043_
timestamp 1644511149
transform -1 0 18216 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _044_
timestamp 1644511149
transform -1 0 3220 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _045_
timestamp 1644511149
transform 1 0 19228 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _046_
timestamp 1644511149
transform 1 0 19412 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _047_
timestamp 1644511149
transform 1 0 18400 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _048_
timestamp 1644511149
transform 1 0 27324 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _049_
timestamp 1644511149
transform -1 0 30176 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _050_
timestamp 1644511149
transform 1 0 16652 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _051_
timestamp 1644511149
transform 1 0 33948 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _052_
timestamp 1644511149
transform 1 0 12880 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _053_
timestamp 1644511149
transform -1 0 18768 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _054_
timestamp 1644511149
transform -1 0 18676 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _055_
timestamp 1644511149
transform 1 0 17848 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _056_
timestamp 1644511149
transform -1 0 6900 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _057_
timestamp 1644511149
transform 1 0 14168 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _058_
timestamp 1644511149
transform -1 0 33856 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _059_
timestamp 1644511149
transform 1 0 17388 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _060_
timestamp 1644511149
transform 1 0 20608 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _061_
timestamp 1644511149
transform -1 0 34316 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _062_
timestamp 1644511149
transform -1 0 3772 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _063_
timestamp 1644511149
transform -1 0 32660 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _064_
timestamp 1644511149
transform -1 0 18216 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _065_
timestamp 1644511149
transform -1 0 11868 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _066_
timestamp 1644511149
transform -1 0 33856 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _067_
timestamp 1644511149
transform 1 0 19412 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _068_
timestamp 1644511149
transform 1 0 17756 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _069_
timestamp 1644511149
transform 1 0 31096 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _070_
timestamp 1644511149
transform 1 0 19964 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _071_
timestamp 1644511149
transform 1 0 17756 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _072_
timestamp 1644511149
transform -1 0 18216 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _073_
timestamp 1644511149
transform 1 0 5428 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _074_
timestamp 1644511149
transform 1 0 17296 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _075_
timestamp 1644511149
transform -1 0 18124 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _076_
timestamp 1644511149
transform -1 0 18768 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _077_
timestamp 1644511149
transform 1 0 24380 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _078_
timestamp 1644511149
transform 1 0 29716 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _079_
timestamp 1644511149
transform 1 0 16928 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _080_
timestamp 1644511149
transform 1 0 18308 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _081_
timestamp 1644511149
transform -1 0 18768 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _082_
timestamp 1644511149
transform 1 0 33948 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _083_
timestamp 1644511149
transform 1 0 17296 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _084_
timestamp 1644511149
transform 1 0 17756 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _085_
timestamp 1644511149
transform -1 0 22172 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _086_
timestamp 1644511149
transform 1 0 17296 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _087_
timestamp 1644511149
transform 1 0 2484 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _088_
timestamp 1644511149
transform -1 0 31188 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _089_
timestamp 1644511149
transform -1 0 33856 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _090_
timestamp 1644511149
transform 1 0 18400 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _091_
timestamp 1644511149
transform 1 0 18400 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _092_
timestamp 1644511149
transform 1 0 6072 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _093_
timestamp 1644511149
transform -1 0 18124 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _094_
timestamp 1644511149
transform -1 0 23552 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _095_
timestamp 1644511149
transform 1 0 1656 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _096_
timestamp 1644511149
transform -1 0 18216 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _097_
timestamp 1644511149
transform 1 0 2392 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _098_
timestamp 1644511149
transform -1 0 17020 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _099_
timestamp 1644511149
transform 1 0 2208 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _100_
timestamp 1644511149
transform 1 0 18952 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _101_
timestamp 1644511149
transform 1 0 1656 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _102_
timestamp 1644511149
transform 1 0 27692 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _103_
timestamp 1644511149
transform -1 0 15640 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _104_
timestamp 1644511149
transform -1 0 16928 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _105_
timestamp 1644511149
transform 1 0 18400 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _106_
timestamp 1644511149
transform -1 0 16008 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _107_
timestamp 1644511149
transform 1 0 10948 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _108_
timestamp 1644511149
transform -1 0 30084 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input1
timestamp 1644511149
transform 1 0 1380 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1644511149
transform 1 0 23276 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1644511149
transform -1 0 11960 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input4 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 34408 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1644511149
transform -1 0 1656 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input6
timestamp 1644511149
transform -1 0 16376 0 -1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input7
timestamp 1644511149
transform 1 0 3772 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input8
timestamp 1644511149
transform -1 0 34408 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input9
timestamp 1644511149
transform 1 0 4876 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1644511149
transform 1 0 34132 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1644511149
transform 1 0 31556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1644511149
transform -1 0 1656 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1644511149
transform 1 0 34132 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input14
timestamp 1644511149
transform -1 0 18952 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input15
timestamp 1644511149
transform -1 0 11224 0 -1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input16
timestamp 1644511149
transform 1 0 30360 0 -1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input17
timestamp 1644511149
transform -1 0 34408 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input18
timestamp 1644511149
transform -1 0 34408 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input19
timestamp 1644511149
transform 1 0 2668 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1644511149
transform 1 0 34132 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input21
timestamp 1644511149
transform -1 0 32660 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input22
timestamp 1644511149
transform 1 0 5704 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input23
timestamp 1644511149
transform -1 0 34408 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1644511149
transform -1 0 16376 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1644511149
transform -1 0 2116 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1644511149
transform -1 0 28704 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1644511149
transform 1 0 34132 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1644511149
transform -1 0 11224 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input29
timestamp 1644511149
transform -1 0 2300 0 -1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1644511149
transform 1 0 9108 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input31
timestamp 1644511149
transform 1 0 31004 0 1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1644511149
transform 1 0 34132 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input33
timestamp 1644511149
transform 1 0 1380 0 -1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input34
timestamp 1644511149
transform 1 0 24380 0 -1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input35
timestamp 1644511149
transform -1 0 34408 0 -1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1644511149
transform -1 0 1656 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input37
timestamp 1644511149
transform -1 0 2300 0 -1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1644511149
transform -1 0 1656 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1644511149
transform 1 0 28612 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1644511149
transform 1 0 1932 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1644511149
transform 1 0 33028 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1644511149
transform -1 0 11316 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input43
timestamp 1644511149
transform -1 0 2300 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input44
timestamp 1644511149
transform 1 0 2484 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input45
timestamp 1644511149
transform 1 0 26956 0 -1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input46
timestamp 1644511149
transform -1 0 33304 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1644511149
transform 1 0 13616 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input48
timestamp 1644511149
transform 1 0 33488 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1644511149
transform 1 0 29716 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1644511149
transform 1 0 21988 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1644511149
transform 1 0 34132 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input52
timestamp 1644511149
transform 1 0 1564 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input53
timestamp 1644511149
transform 1 0 1564 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 1644511149
transform -1 0 22080 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input55
timestamp 1644511149
transform 1 0 29532 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input56
timestamp 1644511149
transform 1 0 33488 0 -1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input57
timestamp 1644511149
transform -1 0 13800 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input58
timestamp 1644511149
transform 1 0 1380 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input59
timestamp 1644511149
transform -1 0 34408 0 1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input60
timestamp 1644511149
transform 1 0 1564 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input61
timestamp 1644511149
transform -1 0 34408 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input62
timestamp 1644511149
transform 1 0 9108 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input63
timestamp 1644511149
transform 1 0 33488 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input64
timestamp 1644511149
transform -1 0 34408 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input65
timestamp 1644511149
transform 1 0 4600 0 -1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input66
timestamp 1644511149
transform -1 0 34408 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input67
timestamp 1644511149
transform 1 0 19228 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input68
timestamp 1644511149
transform -1 0 8096 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input69
timestamp 1644511149
transform -1 0 14904 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input70
timestamp 1644511149
transform 1 0 26956 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input71
timestamp 1644511149
transform 1 0 33488 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input72
timestamp 1644511149
transform -1 0 33304 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input73
timestamp 1644511149
transform 1 0 34132 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input74
timestamp 1644511149
transform 1 0 14904 0 1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input75
timestamp 1644511149
transform 1 0 20608 0 -1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input76
timestamp 1644511149
transform 1 0 19412 0 -1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input77
timestamp 1644511149
transform 1 0 1380 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input78
timestamp 1644511149
transform 1 0 6348 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input79
timestamp 1644511149
transform -1 0 34408 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input80
timestamp 1644511149
transform 1 0 14904 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input81
timestamp 1644511149
transform 1 0 34132 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input82
timestamp 1644511149
transform 1 0 7820 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input83
timestamp 1644511149
transform 1 0 23276 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input84
timestamp 1644511149
transform 1 0 2116 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input85
timestamp 1644511149
transform 1 0 34132 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input86
timestamp 1644511149
transform -1 0 2300 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input87
timestamp 1644511149
transform 1 0 9108 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input88
timestamp 1644511149
transform -1 0 34408 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  output89
timestamp 1644511149
transform 1 0 34040 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp 1644511149
transform 1 0 34040 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output91
timestamp 1644511149
transform -1 0 2852 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output92
timestamp 1644511149
transform -1 0 23000 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output93
timestamp 1644511149
transform -1 0 18492 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output94
timestamp 1644511149
transform -1 0 1748 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output95
timestamp 1644511149
transform -1 0 1748 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output96
timestamp 1644511149
transform -1 0 1748 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output97
timestamp 1644511149
transform -1 0 1748 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output98
timestamp 1644511149
transform 1 0 19228 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output99
timestamp 1644511149
transform 1 0 33488 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output100
timestamp 1644511149
transform 1 0 10212 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output101
timestamp 1644511149
transform 1 0 32292 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output102
timestamp 1644511149
transform 1 0 29716 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output103
timestamp 1644511149
transform -1 0 27508 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output104
timestamp 1644511149
transform -1 0 17020 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output105
timestamp 1644511149
transform 1 0 34040 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output106
timestamp 1644511149
transform -1 0 1748 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output107
timestamp 1644511149
transform -1 0 3404 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output108
timestamp 1644511149
transform -1 0 1748 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output109
timestamp 1644511149
transform 1 0 32936 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output110
timestamp 1644511149
transform 1 0 6532 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output111
timestamp 1644511149
transform -1 0 14444 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output112
timestamp 1644511149
transform -1 0 12052 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output113
timestamp 1644511149
transform 1 0 34040 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output114
timestamp 1644511149
transform -1 0 27508 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output115
timestamp 1644511149
transform -1 0 1748 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output116
timestamp 1644511149
transform 1 0 34040 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output117
timestamp 1644511149
transform 1 0 34040 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output118
timestamp 1644511149
transform 1 0 28060 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output119
timestamp 1644511149
transform 1 0 34040 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output120
timestamp 1644511149
transform -1 0 1748 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output121
timestamp 1644511149
transform -1 0 10120 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output122
timestamp 1644511149
transform 1 0 32384 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output123
timestamp 1644511149
transform -1 0 19780 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output124
timestamp 1644511149
transform 1 0 34040 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output125
timestamp 1644511149
transform -1 0 1748 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output126
timestamp 1644511149
transform 1 0 8280 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output127
timestamp 1644511149
transform 1 0 34040 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output128
timestamp 1644511149
transform 1 0 24380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output129
timestamp 1644511149
transform 1 0 34040 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output130
timestamp 1644511149
transform -1 0 3404 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output131
timestamp 1644511149
transform -1 0 31004 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output132
timestamp 1644511149
transform -1 0 4324 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output133
timestamp 1644511149
transform 1 0 14260 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output134
timestamp 1644511149
transform 1 0 34040 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output135
timestamp 1644511149
transform 1 0 32936 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output136
timestamp 1644511149
transform 1 0 34040 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output137
timestamp 1644511149
transform 1 0 32292 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output138
timestamp 1644511149
transform -1 0 1748 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output139
timestamp 1644511149
transform 1 0 34040 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output140
timestamp 1644511149
transform -1 0 1748 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output141
timestamp 1644511149
transform 1 0 34040 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output142
timestamp 1644511149
transform 1 0 34040 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output143
timestamp 1644511149
transform 1 0 33488 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output144
timestamp 1644511149
transform 1 0 33488 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output145
timestamp 1644511149
transform -1 0 1748 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output146
timestamp 1644511149
transform -1 0 1748 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output147
timestamp 1644511149
transform -1 0 22172 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output148
timestamp 1644511149
transform 1 0 1932 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output149
timestamp 1644511149
transform 1 0 25208 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output150
timestamp 1644511149
transform -1 0 1748 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output151
timestamp 1644511149
transform 1 0 3956 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output152
timestamp 1644511149
transform -1 0 17204 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output153
timestamp 1644511149
transform -1 0 1748 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output154
timestamp 1644511149
transform -1 0 6900 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output155
timestamp 1644511149
transform 1 0 2484 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output156
timestamp 1644511149
transform -1 0 24932 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output157
timestamp 1644511149
transform 1 0 16192 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output158
timestamp 1644511149
transform 1 0 17480 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output159
timestamp 1644511149
transform 1 0 28888 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output160
timestamp 1644511149
transform 1 0 34040 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output161
timestamp 1644511149
transform -1 0 1748 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output162
timestamp 1644511149
transform -1 0 1748 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output163
timestamp 1644511149
transform -1 0 7820 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output164
timestamp 1644511149
transform -1 0 12696 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output165
timestamp 1644511149
transform -1 0 1748 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output166
timestamp 1644511149
transform 1 0 34040 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output167
timestamp 1644511149
transform -1 0 20700 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output168
timestamp 1644511149
transform 1 0 25852 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output169
timestamp 1644511149
transform 1 0 25208 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output170
timestamp 1644511149
transform -1 0 2300 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output171
timestamp 1644511149
transform -1 0 6256 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output172
timestamp 1644511149
transform -1 0 24932 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output173
timestamp 1644511149
transform -1 0 1748 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output174
timestamp 1644511149
transform -1 0 1748 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output175
timestamp 1644511149
transform 1 0 34040 0 -1 17408
box -38 -48 406 592
<< labels >>
rlabel metal3 s 0 19048 800 19168 6 io_dbus_addr[0]
port 0 nsew signal input
rlabel metal2 s 23202 0 23258 800 6 io_dbus_addr[10]
port 1 nsew signal input
rlabel metal2 s 11610 35200 11666 36000 6 io_dbus_addr[11]
port 2 nsew signal input
rlabel metal3 s 35200 4768 36000 4888 6 io_dbus_addr[12]
port 3 nsew signal input
rlabel metal3 s 0 25848 800 25968 6 io_dbus_addr[13]
port 4 nsew signal input
rlabel metal2 s 15474 35200 15530 36000 6 io_dbus_addr[14]
port 5 nsew signal input
rlabel metal2 s 3238 0 3294 800 6 io_dbus_addr[15]
port 6 nsew signal input
rlabel metal3 s 35200 10208 36000 10328 6 io_dbus_addr[16]
port 7 nsew signal input
rlabel metal3 s 0 3408 800 3528 6 io_dbus_addr[17]
port 8 nsew signal input
rlabel metal3 s 0 25168 800 25288 6 io_dbus_addr[18]
port 9 nsew signal input
rlabel metal3 s 0 13608 800 13728 6 io_dbus_addr[19]
port 10 nsew signal input
rlabel metal3 s 35200 26528 36000 26648 6 io_dbus_addr[1]
port 11 nsew signal input
rlabel metal3 s 0 33328 800 33448 6 io_dbus_addr[20]
port 12 nsew signal input
rlabel metal3 s 0 20408 800 20528 6 io_dbus_addr[21]
port 13 nsew signal input
rlabel metal3 s 0 8168 800 8288 6 io_dbus_addr[22]
port 14 nsew signal input
rlabel metal3 s 35200 3408 36000 3528 6 io_dbus_addr[23]
port 15 nsew signal input
rlabel metal2 s 12898 35200 12954 36000 6 io_dbus_addr[24]
port 16 nsew signal input
rlabel metal3 s 0 9528 800 9648 6 io_dbus_addr[25]
port 17 nsew signal input
rlabel metal3 s 0 26528 800 26648 6 io_dbus_addr[26]
port 18 nsew signal input
rlabel metal2 s 3238 35200 3294 36000 6 io_dbus_addr[27]
port 19 nsew signal input
rlabel metal2 s 21914 35200 21970 36000 6 io_dbus_addr[28]
port 20 nsew signal input
rlabel metal2 s 34150 0 34206 800 6 io_dbus_addr[29]
port 21 nsew signal input
rlabel metal2 s 4526 0 4582 800 6 io_dbus_addr[2]
port 22 nsew signal input
rlabel metal3 s 0 4088 800 4208 6 io_dbus_addr[30]
port 23 nsew signal input
rlabel metal2 s 19982 35200 20038 36000 6 io_dbus_addr[31]
port 24 nsew signal input
rlabel metal3 s 35200 25848 36000 25968 6 io_dbus_addr[3]
port 25 nsew signal input
rlabel metal2 s 31574 0 31630 800 6 io_dbus_addr[4]
port 26 nsew signal input
rlabel metal3 s 0 2728 800 2848 6 io_dbus_addr[5]
port 27 nsew signal input
rlabel metal3 s 35200 31288 36000 31408 6 io_dbus_addr[6]
port 28 nsew signal input
rlabel metal2 s 18050 0 18106 800 6 io_dbus_addr[7]
port 29 nsew signal input
rlabel metal2 s 10322 35200 10378 36000 6 io_dbus_addr[8]
port 30 nsew signal input
rlabel metal2 s 30286 35200 30342 36000 6 io_dbus_addr[9]
port 31 nsew signal input
rlabel metal3 s 35200 23808 36000 23928 6 io_dbus_ld_type[0]
port 32 nsew signal input
rlabel metal3 s 35200 34688 36000 34808 6 io_dbus_ld_type[1]
port 33 nsew signal input
rlabel metal2 s 2594 35200 2650 36000 6 io_dbus_ld_type[2]
port 34 nsew signal input
rlabel metal3 s 35200 18368 36000 18488 6 io_dbus_rd_en
port 35 nsew signal input
rlabel metal3 s 35200 31968 36000 32088 6 io_dbus_rdata[0]
port 36 nsew signal tristate
rlabel metal3 s 35200 11568 36000 11688 6 io_dbus_rdata[10]
port 37 nsew signal tristate
rlabel metal3 s 0 34688 800 34808 6 io_dbus_rdata[11]
port 38 nsew signal tristate
rlabel metal2 s 22558 0 22614 800 6 io_dbus_rdata[12]
port 39 nsew signal tristate
rlabel metal2 s 18050 35200 18106 36000 6 io_dbus_rdata[13]
port 40 nsew signal tristate
rlabel metal3 s 0 23128 800 23248 6 io_dbus_rdata[14]
port 41 nsew signal tristate
rlabel metal3 s 0 24488 800 24608 6 io_dbus_rdata[15]
port 42 nsew signal tristate
rlabel metal3 s 0 12248 800 12368 6 io_dbus_rdata[16]
port 43 nsew signal tristate
rlabel metal3 s 0 6128 800 6248 6 io_dbus_rdata[17]
port 44 nsew signal tristate
rlabel metal2 s 18694 35200 18750 36000 6 io_dbus_rdata[18]
port 45 nsew signal tristate
rlabel metal3 s 35200 34008 36000 34128 6 io_dbus_rdata[19]
port 46 nsew signal tristate
rlabel metal2 s 9678 0 9734 800 6 io_dbus_rdata[1]
port 47 nsew signal tristate
rlabel metal2 s 32218 35200 32274 36000 6 io_dbus_rdata[20]
port 48 nsew signal tristate
rlabel metal2 s 29642 35200 29698 36000 6 io_dbus_rdata[21]
port 49 nsew signal tristate
rlabel metal2 s 27066 35200 27122 36000 6 io_dbus_rdata[22]
port 50 nsew signal tristate
rlabel metal2 s 16118 0 16174 800 6 io_dbus_rdata[23]
port 51 nsew signal tristate
rlabel metal3 s 35200 14968 36000 15088 6 io_dbus_rdata[24]
port 52 nsew signal tristate
rlabel metal3 s 0 17688 800 17808 6 io_dbus_rdata[25]
port 53 nsew signal tristate
rlabel metal2 s 2594 0 2650 800 6 io_dbus_rdata[26]
port 54 nsew signal tristate
rlabel metal3 s 0 17008 800 17128 6 io_dbus_rdata[27]
port 55 nsew signal tristate
rlabel metal2 s 32862 0 32918 800 6 io_dbus_rdata[28]
port 56 nsew signal tristate
rlabel metal2 s 6458 35200 6514 36000 6 io_dbus_rdata[29]
port 57 nsew signal tristate
rlabel metal2 s 13542 35200 13598 36000 6 io_dbus_rdata[2]
port 58 nsew signal tristate
rlabel metal2 s 11610 0 11666 800 6 io_dbus_rdata[30]
port 59 nsew signal tristate
rlabel metal3 s 35200 27888 36000 28008 6 io_dbus_rdata[31]
port 60 nsew signal tristate
rlabel metal2 s 27066 0 27122 800 6 io_dbus_rdata[3]
port 61 nsew signal tristate
rlabel metal3 s 0 31288 800 31408 6 io_dbus_rdata[4]
port 62 nsew signal tristate
rlabel metal3 s 35200 8848 36000 8968 6 io_dbus_rdata[5]
port 63 nsew signal tristate
rlabel metal3 s 35200 17688 36000 17808 6 io_dbus_rdata[6]
port 64 nsew signal tristate
rlabel metal2 s 27710 0 27766 800 6 io_dbus_rdata[7]
port 65 nsew signal tristate
rlabel metal3 s 35200 4088 36000 4208 6 io_dbus_rdata[8]
port 66 nsew signal tristate
rlabel metal3 s 0 14288 800 14408 6 io_dbus_rdata[9]
port 67 nsew signal tristate
rlabel metal2 s 31574 35200 31630 36000 6 io_dbus_st_type[0]
port 68 nsew signal input
rlabel metal2 s 5170 35200 5226 36000 6 io_dbus_st_type[1]
port 69 nsew signal input
rlabel metal2 s 9678 35200 9734 36000 6 io_dbus_valid
port 70 nsew signal tristate
rlabel metal3 s 35200 8168 36000 8288 6 io_dbus_wdata[0]
port 71 nsew signal input
rlabel metal2 s 16762 0 16818 800 6 io_dbus_wdata[10]
port 72 nsew signal input
rlabel metal3 s 0 688 800 808 6 io_dbus_wdata[11]
port 73 nsew signal input
rlabel metal2 s 28354 35200 28410 36000 6 io_dbus_wdata[12]
port 74 nsew signal input
rlabel metal3 s 35200 29248 36000 29368 6 io_dbus_wdata[13]
port 75 nsew signal input
rlabel metal2 s 10966 0 11022 800 6 io_dbus_wdata[14]
port 76 nsew signal input
rlabel metal3 s 0 29928 800 30048 6 io_dbus_wdata[15]
port 77 nsew signal input
rlabel metal2 s 9034 35200 9090 36000 6 io_dbus_wdata[16]
port 78 nsew signal input
rlabel metal2 s 30930 35200 30986 36000 6 io_dbus_wdata[17]
port 79 nsew signal input
rlabel metal3 s 35200 19048 36000 19168 6 io_dbus_wdata[18]
port 80 nsew signal input
rlabel metal3 s 0 31968 800 32088 6 io_dbus_wdata[19]
port 81 nsew signal input
rlabel metal2 s 23846 35200 23902 36000 6 io_dbus_wdata[1]
port 82 nsew signal input
rlabel metal3 s 35200 21088 36000 21208 6 io_dbus_wdata[20]
port 83 nsew signal input
rlabel metal3 s 0 14968 800 15088 6 io_dbus_wdata[21]
port 84 nsew signal input
rlabel metal2 s 662 35200 718 36000 6 io_dbus_wdata[22]
port 85 nsew signal input
rlabel metal3 s 0 10208 800 10328 6 io_dbus_wdata[23]
port 86 nsew signal input
rlabel metal2 s 28354 0 28410 800 6 io_dbus_wdata[24]
port 87 nsew signal input
rlabel metal3 s 0 18368 800 18488 6 io_dbus_wdata[25]
port 88 nsew signal input
rlabel metal2 s 33506 35200 33562 36000 6 io_dbus_wdata[26]
port 89 nsew signal input
rlabel metal2 s 10966 35200 11022 36000 6 io_dbus_wdata[27]
port 90 nsew signal input
rlabel metal2 s 1306 0 1362 800 6 io_dbus_wdata[28]
port 91 nsew signal input
rlabel metal3 s 0 2048 800 2168 6 io_dbus_wdata[29]
port 92 nsew signal input
rlabel metal2 s 26422 35200 26478 36000 6 io_dbus_wdata[2]
port 93 nsew signal input
rlabel metal3 s 35200 1368 36000 1488 6 io_dbus_wdata[30]
port 94 nsew signal input
rlabel metal2 s 13542 0 13598 800 6 io_dbus_wdata[31]
port 95 nsew signal input
rlabel metal3 s 35200 688 36000 808 6 io_dbus_wdata[3]
port 96 nsew signal input
rlabel metal2 s 29642 0 29698 800 6 io_dbus_wdata[4]
port 97 nsew signal input
rlabel metal2 s 21914 0 21970 800 6 io_dbus_wdata[5]
port 98 nsew signal input
rlabel metal3 s 35200 19728 36000 19848 6 io_dbus_wdata[6]
port 99 nsew signal input
rlabel metal3 s 0 28568 800 28688 6 io_dbus_wdata[7]
port 100 nsew signal input
rlabel metal3 s 0 12928 800 13048 6 io_dbus_wdata[8]
port 101 nsew signal input
rlabel metal2 s 21270 35200 21326 36000 6 io_dbus_wdata[9]
port 102 nsew signal input
rlabel metal2 s 28998 0 29054 800 6 io_dbus_wr_en
port 103 nsew signal input
rlabel metal3 s 35200 35368 36000 35488 6 io_wbm_ack_i
port 104 nsew signal input
rlabel metal2 s 12898 0 12954 800 6 io_wbm_data_i[0]
port 105 nsew signal input
rlabel metal3 s 0 11568 800 11688 6 io_wbm_data_i[10]
port 106 nsew signal input
rlabel metal3 s 35200 30608 36000 30728 6 io_wbm_data_i[11]
port 107 nsew signal input
rlabel metal2 s 18 35200 74 36000 6 io_wbm_data_i[12]
port 108 nsew signal input
rlabel metal3 s 35200 13608 36000 13728 6 io_wbm_data_i[13]
port 109 nsew signal input
rlabel metal2 s 9034 0 9090 800 6 io_wbm_data_i[14]
port 110 nsew signal input
rlabel metal3 s 35200 20408 36000 20528 6 io_wbm_data_i[15]
port 111 nsew signal input
rlabel metal2 s 35438 0 35494 800 6 io_wbm_data_i[16]
port 112 nsew signal input
rlabel metal2 s 4526 35200 4582 36000 6 io_wbm_data_i[17]
port 113 nsew signal input
rlabel metal3 s 35200 22448 36000 22568 6 io_wbm_data_i[18]
port 114 nsew signal input
rlabel metal2 s 18694 0 18750 800 6 io_wbm_data_i[19]
port 115 nsew signal input
rlabel metal2 s 7746 0 7802 800 6 io_wbm_data_i[1]
port 116 nsew signal input
rlabel metal2 s 14186 35200 14242 36000 6 io_wbm_data_i[20]
port 117 nsew signal input
rlabel metal2 s 26422 0 26478 800 6 io_wbm_data_i[21]
port 118 nsew signal input
rlabel metal2 s 33506 0 33562 800 6 io_wbm_data_i[22]
port 119 nsew signal input
rlabel metal2 s 34794 35200 34850 36000 6 io_wbm_data_i[23]
port 120 nsew signal input
rlabel metal3 s 35200 14288 36000 14408 6 io_wbm_data_i[24]
port 121 nsew signal input
rlabel metal2 s 14830 35200 14886 36000 6 io_wbm_data_i[25]
port 122 nsew signal input
rlabel metal2 s 20626 35200 20682 36000 6 io_wbm_data_i[26]
port 123 nsew signal input
rlabel metal2 s 19338 35200 19394 36000 6 io_wbm_data_i[27]
port 124 nsew signal input
rlabel metal3 s 0 19728 800 19848 6 io_wbm_data_i[28]
port 125 nsew signal input
rlabel metal2 s 5814 0 5870 800 6 io_wbm_data_i[29]
port 126 nsew signal input
rlabel metal3 s 35200 6128 36000 6248 6 io_wbm_data_i[2]
port 127 nsew signal input
rlabel metal2 s 14830 0 14886 800 6 io_wbm_data_i[30]
port 128 nsew signal input
rlabel metal3 s 35200 29928 36000 30048 6 io_wbm_data_i[31]
port 129 nsew signal input
rlabel metal2 s 7746 35200 7802 36000 6 io_wbm_data_i[3]
port 130 nsew signal input
rlabel metal2 s 23202 35200 23258 36000 6 io_wbm_data_i[4]
port 131 nsew signal input
rlabel metal3 s 0 34008 800 34128 6 io_wbm_data_i[5]
port 132 nsew signal input
rlabel metal3 s 35200 9528 36000 9648 6 io_wbm_data_i[6]
port 133 nsew signal input
rlabel metal3 s 0 1368 800 1488 6 io_wbm_data_i[7]
port 134 nsew signal input
rlabel metal2 s 8390 35200 8446 36000 6 io_wbm_data_i[8]
port 135 nsew signal input
rlabel metal3 s 35200 15648 36000 15768 6 io_wbm_data_i[9]
port 136 nsew signal input
rlabel metal3 s 35200 2048 36000 2168 6 io_wbm_m2s_addr[0]
port 137 nsew signal tristate
rlabel metal2 s 19338 0 19394 800 6 io_wbm_m2s_addr[10]
port 138 nsew signal tristate
rlabel metal3 s 35200 28568 36000 28688 6 io_wbm_m2s_addr[11]
port 139 nsew signal tristate
rlabel metal3 s 0 4768 800 4888 6 io_wbm_m2s_addr[12]
port 140 nsew signal tristate
rlabel metal2 s 8390 0 8446 800 6 io_wbm_m2s_addr[13]
port 141 nsew signal tristate
rlabel metal3 s 35200 12248 36000 12368 6 io_wbm_m2s_addr[14]
port 142 nsew signal tristate
rlabel metal2 s 23846 0 23902 800 6 io_wbm_m2s_addr[15]
port 143 nsew signal tristate
rlabel metal3 s 35200 2728 36000 2848 6 io_wbm_m2s_addr[1]
port 144 nsew signal tristate
rlabel metal2 s 1306 35200 1362 36000 6 io_wbm_m2s_addr[2]
port 145 nsew signal tristate
rlabel metal2 s 30286 0 30342 800 6 io_wbm_m2s_addr[3]
port 146 nsew signal tristate
rlabel metal2 s 3882 0 3938 800 6 io_wbm_m2s_addr[4]
port 147 nsew signal tristate
rlabel metal2 s 14186 0 14242 800 6 io_wbm_m2s_addr[5]
port 148 nsew signal tristate
rlabel metal3 s 35200 7488 36000 7608 6 io_wbm_m2s_addr[6]
port 149 nsew signal tristate
rlabel metal3 s 35200 33328 36000 33448 6 io_wbm_m2s_addr[7]
port 150 nsew signal tristate
rlabel metal3 s 35200 23128 36000 23248 6 io_wbm_m2s_addr[8]
port 151 nsew signal tristate
rlabel metal2 s 32218 0 32274 800 6 io_wbm_m2s_addr[9]
port 152 nsew signal tristate
rlabel metal3 s 0 15648 800 15768 6 io_wbm_m2s_data[0]
port 153 nsew signal tristate
rlabel metal3 s 35200 12928 36000 13048 6 io_wbm_m2s_data[10]
port 154 nsew signal tristate
rlabel metal2 s 662 0 718 800 6 io_wbm_m2s_data[11]
port 155 nsew signal tristate
rlabel metal3 s 35200 25168 36000 25288 6 io_wbm_m2s_data[12]
port 156 nsew signal tristate
rlabel metal2 s 35438 35200 35494 36000 6 io_wbm_m2s_data[13]
port 157 nsew signal tristate
rlabel metal2 s 34794 0 34850 800 6 io_wbm_m2s_data[14]
port 158 nsew signal tristate
rlabel metal2 s 34150 35200 34206 36000 6 io_wbm_m2s_data[15]
port 159 nsew signal tristate
rlabel metal3 s 0 22448 800 22568 6 io_wbm_m2s_data[16]
port 160 nsew signal tristate
rlabel metal3 s 0 23808 800 23928 6 io_wbm_m2s_data[17]
port 161 nsew signal tristate
rlabel metal2 s 21270 0 21326 800 6 io_wbm_m2s_data[18]
port 162 nsew signal tristate
rlabel metal2 s 18 0 74 800 6 io_wbm_m2s_data[19]
port 163 nsew signal tristate
rlabel metal2 s 25134 0 25190 800 6 io_wbm_m2s_data[1]
port 164 nsew signal tristate
rlabel metal3 s 0 27888 800 28008 6 io_wbm_m2s_data[20]
port 165 nsew signal tristate
rlabel metal2 s 3882 35200 3938 36000 6 io_wbm_m2s_data[21]
port 166 nsew signal tristate
rlabel metal2 s 16762 35200 16818 36000 6 io_wbm_m2s_data[22]
port 167 nsew signal tristate
rlabel metal3 s 0 21088 800 21208 6 io_wbm_m2s_data[23]
port 168 nsew signal tristate
rlabel metal2 s 6458 0 6514 800 6 io_wbm_m2s_data[24]
port 169 nsew signal tristate
rlabel metal2 s 1950 0 2006 800 6 io_wbm_m2s_data[25]
port 170 nsew signal tristate
rlabel metal2 s 24490 35200 24546 36000 6 io_wbm_m2s_data[26]
port 171 nsew signal tristate
rlabel metal2 s 16118 35200 16174 36000 6 io_wbm_m2s_data[27]
port 172 nsew signal tristate
rlabel metal2 s 17406 0 17462 800 6 io_wbm_m2s_data[28]
port 173 nsew signal tristate
rlabel metal2 s 28998 35200 29054 36000 6 io_wbm_m2s_data[29]
port 174 nsew signal tristate
rlabel metal3 s 35200 6808 36000 6928 6 io_wbm_m2s_data[2]
port 175 nsew signal tristate
rlabel metal3 s 0 29248 800 29368 6 io_wbm_m2s_data[30]
port 176 nsew signal tristate
rlabel metal3 s 0 7488 800 7608 6 io_wbm_m2s_data[31]
port 177 nsew signal tristate
rlabel metal2 s 7102 0 7158 800 6 io_wbm_m2s_data[3]
port 178 nsew signal tristate
rlabel metal2 s 12254 0 12310 800 6 io_wbm_m2s_data[4]
port 179 nsew signal tristate
rlabel metal3 s 0 6808 800 6928 6 io_wbm_m2s_data[5]
port 180 nsew signal tristate
rlabel metal3 s 35200 24488 36000 24608 6 io_wbm_m2s_data[6]
port 181 nsew signal tristate
rlabel metal2 s 19982 0 20038 800 6 io_wbm_m2s_data[7]
port 182 nsew signal tristate
rlabel metal2 s 25778 35200 25834 36000 6 io_wbm_m2s_data[8]
port 183 nsew signal tristate
rlabel metal2 s 25134 35200 25190 36000 6 io_wbm_m2s_data[9]
port 184 nsew signal tristate
rlabel metal3 s 0 35368 800 35488 6 io_wbm_m2s_sel[0]
port 185 nsew signal tristate
rlabel metal2 s 5814 35200 5870 36000 6 io_wbm_m2s_sel[1]
port 186 nsew signal tristate
rlabel metal2 s 24490 0 24546 800 6 io_wbm_m2s_sel[2]
port 187 nsew signal tristate
rlabel metal3 s 0 8848 800 8968 6 io_wbm_m2s_sel[3]
port 188 nsew signal tristate
rlabel metal3 s 0 30608 800 30728 6 io_wbm_m2s_stb
port 189 nsew signal tristate
rlabel metal3 s 35200 17008 36000 17128 6 io_wbm_m2s_we
port 190 nsew signal tristate
rlabel metal4 s 6576 2128 6896 33776 6 vccd1
port 191 nsew power input
rlabel metal4 s 17840 2128 18160 33776 6 vccd1
port 191 nsew power input
rlabel metal4 s 29104 2128 29424 33776 6 vccd1
port 191 nsew power input
rlabel metal4 s 12208 2128 12528 33776 6 vssd1
port 192 nsew ground input
rlabel metal4 s 23472 2128 23792 33776 6 vssd1
port 192 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 36000 36000
<< end >>
