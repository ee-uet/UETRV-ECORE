magic
tech sky130A
magscale 1 2
timestamp 1647505415
<< viali >>
rect 2421 27557 2455 27591
rect 3985 27557 4019 27591
rect 16773 27557 16807 27591
rect 19441 27557 19475 27591
rect 21833 27557 21867 27591
rect 22385 27557 22419 27591
rect 23949 27557 23983 27591
rect 25513 27557 25547 27591
rect 25881 27557 25915 27591
rect 27813 27557 27847 27591
rect 28273 27557 28307 27591
rect 1685 27421 1719 27455
rect 2789 27421 2823 27455
rect 10517 27421 10551 27455
rect 10977 27421 11011 27455
rect 16957 27421 16991 27455
rect 22753 27421 22787 27455
rect 24685 27421 24719 27455
rect 25329 27421 25363 27455
rect 28089 27421 28123 27455
rect 3157 27353 3191 27387
rect 10701 27353 10735 27387
rect 25053 27353 25087 27387
rect 1777 27285 1811 27319
rect 22845 27285 22879 27319
rect 2329 27081 2363 27115
rect 23489 27081 23523 27115
rect 25145 27081 25179 27115
rect 28273 27081 28307 27115
rect 1409 26945 1443 26979
rect 1961 26945 1995 26979
rect 22376 26945 22410 26979
rect 23765 26945 23799 26979
rect 24032 26945 24066 26979
rect 28089 26945 28123 26979
rect 22109 26877 22143 26911
rect 1593 26741 1627 26775
rect 28365 26537 28399 26571
rect 1409 26333 1443 26367
rect 27813 25245 27847 25279
rect 28365 25245 28399 25279
rect 28181 25109 28215 25143
rect 1409 24769 1443 24803
rect 1961 24769 1995 24803
rect 14933 24769 14967 24803
rect 1593 24565 1627 24599
rect 14749 24565 14783 24599
rect 14381 24157 14415 24191
rect 14648 24157 14682 24191
rect 16681 24157 16715 24191
rect 15761 24021 15795 24055
rect 16129 24021 16163 24055
rect 16865 24021 16899 24055
rect 17233 24021 17267 24055
rect 14657 23817 14691 23851
rect 16313 23817 16347 23851
rect 15301 23749 15335 23783
rect 20913 23749 20947 23783
rect 14473 23681 14507 23715
rect 15393 23681 15427 23715
rect 16129 23681 16163 23715
rect 16948 23681 16982 23715
rect 19533 23681 19567 23715
rect 20729 23681 20763 23715
rect 14289 23613 14323 23647
rect 15485 23613 15519 23647
rect 15945 23613 15979 23647
rect 16681 23613 16715 23647
rect 14933 23545 14967 23579
rect 19349 23545 19383 23579
rect 1409 23477 1443 23511
rect 18061 23477 18095 23511
rect 19993 23477 20027 23511
rect 28365 23477 28399 23511
rect 15301 23273 15335 23307
rect 16221 23273 16255 23307
rect 15577 23137 15611 23171
rect 16773 23137 16807 23171
rect 12817 23069 12851 23103
rect 13461 23069 13495 23103
rect 15761 23069 15795 23103
rect 16589 23069 16623 23103
rect 17785 23069 17819 23103
rect 18429 23069 18463 23103
rect 18889 23069 18923 23103
rect 20085 23069 20119 23103
rect 20269 23069 20303 23103
rect 15945 23001 15979 23035
rect 17417 23001 17451 23035
rect 19533 23001 19567 23035
rect 19717 23001 19751 23035
rect 13001 22933 13035 22967
rect 13277 22933 13311 22967
rect 16681 22933 16715 22967
rect 17325 22933 17359 22967
rect 17969 22933 18003 22967
rect 18245 22933 18279 22967
rect 18705 22933 18739 22967
rect 20453 22933 20487 22967
rect 12633 22729 12667 22763
rect 14289 22729 14323 22763
rect 15025 22729 15059 22763
rect 16129 22729 16163 22763
rect 13154 22661 13188 22695
rect 14933 22661 14967 22695
rect 15761 22661 15795 22695
rect 18604 22661 18638 22695
rect 12357 22593 12391 22627
rect 12449 22593 12483 22627
rect 12909 22593 12943 22627
rect 15577 22593 15611 22627
rect 15853 22593 15887 22627
rect 15945 22593 15979 22627
rect 17805 22593 17839 22627
rect 18061 22593 18095 22627
rect 18337 22593 18371 22627
rect 21209 22593 21243 22627
rect 21465 22593 21499 22627
rect 15117 22525 15151 22559
rect 20085 22457 20119 22491
rect 10517 22389 10551 22423
rect 14565 22389 14599 22423
rect 16681 22389 16715 22423
rect 19717 22389 19751 22423
rect 16221 22185 16255 22219
rect 18889 22185 18923 22219
rect 20269 22185 20303 22219
rect 21281 22185 21315 22219
rect 16773 22049 16807 22083
rect 19901 22049 19935 22083
rect 20729 22049 20763 22083
rect 20913 22049 20947 22083
rect 7849 21981 7883 22015
rect 9597 21981 9631 22015
rect 10333 21981 10367 22015
rect 12081 21981 12115 22015
rect 12357 21981 12391 22015
rect 15669 21981 15703 22015
rect 17332 21981 17366 22015
rect 17463 21981 17497 22015
rect 17555 21981 17589 22015
rect 17690 21981 17724 22015
rect 17790 21981 17824 22015
rect 18613 21981 18647 22015
rect 18705 21981 18739 22015
rect 20637 21981 20671 22015
rect 21465 21981 21499 22015
rect 10149 21913 10183 21947
rect 11814 21913 11848 21947
rect 12624 21913 12658 21947
rect 15424 21913 15458 21947
rect 19717 21913 19751 21947
rect 8033 21845 8067 21879
rect 9413 21845 9447 21879
rect 10701 21845 10735 21879
rect 13737 21845 13771 21879
rect 14289 21845 14323 21879
rect 16589 21845 16623 21879
rect 16681 21845 16715 21879
rect 17969 21845 18003 21879
rect 19257 21845 19291 21879
rect 19625 21845 19659 21879
rect 21741 21845 21775 21879
rect 10701 21641 10735 21675
rect 11989 21641 12023 21675
rect 12909 21641 12943 21675
rect 14013 21641 14047 21675
rect 16681 21641 16715 21675
rect 19165 21641 19199 21675
rect 21373 21641 21407 21675
rect 9566 21573 9600 21607
rect 11897 21573 11931 21607
rect 15117 21573 15151 21607
rect 17776 21573 17810 21607
rect 7665 21505 7699 21539
rect 7932 21505 7966 21539
rect 10977 21505 11011 21539
rect 12725 21505 12759 21539
rect 13921 21505 13955 21539
rect 15025 21505 15059 21539
rect 15945 21505 15979 21539
rect 16129 21505 16163 21539
rect 16865 21505 16899 21539
rect 17509 21505 17543 21539
rect 19349 21505 19383 21539
rect 19533 21505 19567 21539
rect 19993 21505 20027 21539
rect 20177 21505 20211 21539
rect 20913 21505 20947 21539
rect 9321 21437 9355 21471
rect 12173 21437 12207 21471
rect 12541 21437 12575 21471
rect 14197 21437 14231 21471
rect 14933 21437 14967 21471
rect 15761 21437 15795 21471
rect 13553 21369 13587 21403
rect 15485 21369 15519 21403
rect 1409 21301 1443 21335
rect 9045 21301 9079 21335
rect 11161 21301 11195 21335
rect 11529 21301 11563 21335
rect 13277 21301 13311 21335
rect 17233 21301 17267 21335
rect 18889 21301 18923 21335
rect 20361 21301 20395 21335
rect 21097 21301 21131 21335
rect 7573 21097 7607 21131
rect 11621 21097 11655 21131
rect 18889 21097 18923 21131
rect 19717 21097 19751 21131
rect 24041 21097 24075 21131
rect 7849 21029 7883 21063
rect 10425 21029 10459 21063
rect 15853 21029 15887 21063
rect 16865 21029 16899 21063
rect 19993 21029 20027 21063
rect 6929 20961 6963 20995
rect 7205 20961 7239 20995
rect 8493 20961 8527 20995
rect 9965 20961 9999 20995
rect 15025 20961 15059 20995
rect 16313 20961 16347 20995
rect 17509 20961 17543 20995
rect 18245 20961 18279 20995
rect 18429 20961 18463 20995
rect 19349 20961 19383 20995
rect 20545 20961 20579 20995
rect 7389 20893 7423 20927
rect 8309 20893 8343 20927
rect 9781 20893 9815 20927
rect 10885 20893 10919 20927
rect 10977 20893 11011 20927
rect 11161 20893 11195 20927
rect 11437 20893 11471 20927
rect 11897 20893 11931 20927
rect 15301 20893 15335 20927
rect 15669 20893 15703 20927
rect 17325 20893 17359 20927
rect 19533 20893 19567 20927
rect 22118 20893 22152 20927
rect 22385 20893 22419 20927
rect 22661 20893 22695 20927
rect 9873 20825 9907 20859
rect 12142 20825 12176 20859
rect 17141 20825 17175 20859
rect 22906 20825 22940 20859
rect 8217 20757 8251 20791
rect 9413 20757 9447 20791
rect 13277 20757 13311 20791
rect 14105 20757 14139 20791
rect 16405 20757 16439 20791
rect 16497 20757 16531 20791
rect 17877 20757 17911 20791
rect 18521 20757 18555 20791
rect 20361 20757 20395 20791
rect 20453 20757 20487 20791
rect 21005 20757 21039 20791
rect 9689 20553 9723 20587
rect 11161 20553 11195 20587
rect 12265 20553 12299 20587
rect 15025 20553 15059 20587
rect 18521 20553 18555 20587
rect 19625 20553 19659 20587
rect 19901 20553 19935 20587
rect 21097 20553 21131 20587
rect 8953 20485 8987 20519
rect 13277 20485 13311 20519
rect 15853 20485 15887 20519
rect 18889 20485 18923 20519
rect 22946 20485 22980 20519
rect 7104 20417 7138 20451
rect 9505 20417 9539 20451
rect 10333 20417 10367 20451
rect 10885 20417 10919 20451
rect 10977 20417 11011 20451
rect 12173 20417 12207 20451
rect 13737 20417 13771 20451
rect 14289 20417 14323 20451
rect 14933 20417 14967 20451
rect 15669 20417 15703 20451
rect 16681 20417 16715 20451
rect 16937 20417 16971 20451
rect 18700 20417 18734 20451
rect 18797 20417 18831 20451
rect 19072 20417 19106 20451
rect 19165 20417 19199 20451
rect 19441 20417 19475 20451
rect 20269 20417 20303 20451
rect 20913 20417 20947 20451
rect 6837 20349 6871 20383
rect 9321 20349 9355 20383
rect 10149 20349 10183 20383
rect 12357 20349 12391 20383
rect 15209 20349 15243 20383
rect 20361 20349 20395 20383
rect 20545 20349 20579 20383
rect 23213 20349 23247 20383
rect 11805 20281 11839 20315
rect 13461 20281 13495 20315
rect 21833 20281 21867 20315
rect 8217 20213 8251 20247
rect 8861 20213 8895 20247
rect 10517 20213 10551 20247
rect 13921 20213 13955 20247
rect 14565 20213 14599 20247
rect 18061 20213 18095 20247
rect 6929 20009 6963 20043
rect 15485 20009 15519 20043
rect 17141 20009 17175 20043
rect 18613 20009 18647 20043
rect 19349 20009 19383 20043
rect 7849 19941 7883 19975
rect 21465 19941 21499 19975
rect 8401 19873 8435 19907
rect 14105 19873 14139 19907
rect 22017 19873 22051 19907
rect 1409 19805 1443 19839
rect 1685 19805 1719 19839
rect 6745 19805 6779 19839
rect 7205 19805 7239 19839
rect 7389 19805 7423 19839
rect 7573 19805 7607 19839
rect 9045 19805 9079 19839
rect 10977 19805 11011 19839
rect 13461 19805 13495 19839
rect 13737 19805 13771 19839
rect 14361 19805 14395 19839
rect 15945 19805 15979 19839
rect 16129 19805 16163 19839
rect 16221 19805 16255 19839
rect 17049 19805 17083 19839
rect 17969 19805 18003 19839
rect 18117 19805 18151 19839
rect 18337 19805 18371 19839
rect 18434 19805 18468 19839
rect 22385 19805 22419 19839
rect 9312 19737 9346 19771
rect 11244 19737 11278 19771
rect 18245 19737 18279 19771
rect 20085 19737 20119 19771
rect 21649 19737 21683 19771
rect 22652 19737 22686 19771
rect 8217 19669 8251 19703
rect 8309 19669 8343 19703
rect 10425 19669 10459 19703
rect 12357 19669 12391 19703
rect 15761 19669 15795 19703
rect 17509 19669 17543 19703
rect 19809 19669 19843 19703
rect 20545 19669 20579 19703
rect 21097 19669 21131 19703
rect 23765 19669 23799 19703
rect 1409 19465 1443 19499
rect 6837 19465 6871 19499
rect 9321 19465 9355 19499
rect 10425 19465 10459 19499
rect 11529 19465 11563 19499
rect 13645 19465 13679 19499
rect 15485 19465 15519 19499
rect 16221 19465 16255 19499
rect 17049 19465 17083 19499
rect 18889 19465 18923 19499
rect 22569 19465 22603 19499
rect 10793 19397 10827 19431
rect 22845 19397 22879 19431
rect 24225 19397 24259 19431
rect 7021 19329 7055 19363
rect 8861 19329 8895 19363
rect 9045 19329 9079 19363
rect 9505 19329 9539 19363
rect 10885 19329 10919 19363
rect 11713 19329 11747 19363
rect 12449 19329 12483 19363
rect 13461 19329 13495 19363
rect 15301 19329 15335 19363
rect 15577 19329 15611 19363
rect 16037 19329 16071 19363
rect 16313 19329 16347 19363
rect 16865 19329 16899 19363
rect 17141 19329 17175 19363
rect 17509 19329 17543 19363
rect 17776 19329 17810 19363
rect 20370 19329 20404 19363
rect 20637 19329 20671 19363
rect 21097 19329 21131 19363
rect 21281 19329 21315 19363
rect 21925 19329 21959 19363
rect 22088 19335 22122 19369
rect 22201 19329 22235 19363
rect 22313 19329 22347 19363
rect 23029 19329 23063 19363
rect 23213 19329 23247 19363
rect 23489 19329 23523 19363
rect 23673 19329 23707 19363
rect 7757 19261 7791 19295
rect 8677 19261 8711 19295
rect 9873 19261 9907 19295
rect 10977 19261 11011 19295
rect 12173 19261 12207 19295
rect 13277 19261 13311 19295
rect 14749 19261 14783 19295
rect 24685 19261 24719 19295
rect 15853 19193 15887 19227
rect 15117 19125 15151 19159
rect 16681 19125 16715 19159
rect 19257 19125 19291 19159
rect 21465 19125 21499 19159
rect 23857 19125 23891 19159
rect 24317 19125 24351 19159
rect 8953 18921 8987 18955
rect 12449 18921 12483 18955
rect 13093 18921 13127 18955
rect 17877 18921 17911 18955
rect 18705 18921 18739 18955
rect 21925 18921 21959 18955
rect 25789 18921 25823 18955
rect 15577 18853 15611 18887
rect 22845 18853 22879 18887
rect 9505 18785 9539 18819
rect 10977 18785 11011 18819
rect 14105 18785 14139 18819
rect 15117 18785 15151 18819
rect 19441 18785 19475 18819
rect 1409 18717 1443 18751
rect 6653 18717 6687 18751
rect 6920 18717 6954 18751
rect 9321 18717 9355 18751
rect 10885 18717 10919 18751
rect 11437 18717 11471 18751
rect 14381 18717 14415 18751
rect 14470 18717 14504 18751
rect 14565 18717 14599 18751
rect 14749 18717 14783 18751
rect 15025 18717 15059 18751
rect 15301 18717 15335 18751
rect 15393 18717 15427 18751
rect 16129 18717 16163 18751
rect 16405 18717 16439 18751
rect 17233 18717 17267 18751
rect 17417 18717 17451 18751
rect 17509 18717 17543 18751
rect 17601 18717 17635 18751
rect 18153 18717 18187 18751
rect 18797 18717 18831 18751
rect 20361 18717 20395 18751
rect 20453 18717 20487 18751
rect 20545 18717 20579 18751
rect 20729 18717 20763 18751
rect 21281 18717 21315 18751
rect 21465 18717 21499 18751
rect 21557 18717 21591 18751
rect 21649 18717 21683 18751
rect 22385 18717 22419 18751
rect 23213 18717 23247 18751
rect 23376 18717 23410 18751
rect 23476 18717 23510 18751
rect 23601 18717 23635 18751
rect 24409 18717 24443 18751
rect 9413 18649 9447 18683
rect 12265 18649 12299 18683
rect 12909 18649 12943 18683
rect 13109 18649 13143 18683
rect 16313 18649 16347 18683
rect 19625 18649 19659 18683
rect 19809 18649 19843 18683
rect 22201 18649 22235 18683
rect 23857 18649 23891 18683
rect 24654 18649 24688 18683
rect 8033 18581 8067 18615
rect 10425 18581 10459 18615
rect 10793 18581 10827 18615
rect 11621 18581 11655 18615
rect 12465 18581 12499 18615
rect 12633 18581 12667 18615
rect 13277 18581 13311 18615
rect 15945 18581 15979 18615
rect 16957 18581 16991 18615
rect 18337 18581 18371 18615
rect 20085 18581 20119 18615
rect 22569 18581 22603 18615
rect 7113 18377 7147 18411
rect 7481 18377 7515 18411
rect 7849 18377 7883 18411
rect 8585 18377 8619 18411
rect 9597 18377 9631 18411
rect 12909 18377 12943 18411
rect 13829 18377 13863 18411
rect 19625 18377 19659 18411
rect 22477 18377 22511 18411
rect 8677 18309 8711 18343
rect 13185 18309 13219 18343
rect 13401 18309 13435 18343
rect 17785 18309 17819 18343
rect 20269 18309 20303 18343
rect 20453 18309 20487 18343
rect 21281 18309 21315 18343
rect 23489 18309 23523 18343
rect 24010 18309 24044 18343
rect 5753 18241 5787 18275
rect 6929 18241 6963 18275
rect 9505 18241 9539 18275
rect 10609 18241 10643 18275
rect 11785 18241 11819 18275
rect 14013 18241 14047 18275
rect 14105 18241 14139 18275
rect 14381 18241 14415 18275
rect 14841 18241 14875 18275
rect 14933 18241 14967 18275
rect 15209 18241 15243 18275
rect 16037 18241 16071 18275
rect 16957 18241 16991 18275
rect 18245 18241 18279 18275
rect 18501 18241 18535 18275
rect 20637 18241 20671 18275
rect 21097 18241 21131 18275
rect 21833 18241 21867 18275
rect 22017 18241 22051 18275
rect 22109 18241 22143 18275
rect 22201 18241 22235 18275
rect 22845 18241 22879 18275
rect 23024 18241 23058 18275
rect 23121 18241 23155 18275
rect 23259 18241 23293 18275
rect 23765 18241 23799 18275
rect 6009 18173 6043 18207
rect 6745 18173 6779 18207
rect 7941 18173 7975 18207
rect 8125 18173 8159 18207
rect 9689 18173 9723 18207
rect 10425 18173 10459 18207
rect 11529 18173 11563 18207
rect 15117 18173 15151 18207
rect 16313 18173 16347 18207
rect 16681 18173 16715 18207
rect 13553 18105 13587 18139
rect 14289 18105 14323 18139
rect 4629 18037 4663 18071
rect 9137 18037 9171 18071
rect 10793 18037 10827 18071
rect 13369 18037 13403 18071
rect 14657 18037 14691 18071
rect 19993 18037 20027 18071
rect 20913 18037 20947 18071
rect 25145 18037 25179 18071
rect 8125 17833 8159 17867
rect 10609 17833 10643 17867
rect 11161 17833 11195 17867
rect 12357 17833 12391 17867
rect 12817 17833 12851 17867
rect 13461 17833 13495 17867
rect 18429 17833 18463 17867
rect 21189 17833 21223 17867
rect 23305 17833 23339 17867
rect 10333 17765 10367 17799
rect 13001 17765 13035 17799
rect 13645 17765 13679 17799
rect 22293 17765 22327 17799
rect 15485 17697 15519 17731
rect 17969 17697 18003 17731
rect 19809 17697 19843 17731
rect 6009 17629 6043 17663
rect 8953 17629 8987 17663
rect 10977 17629 11011 17663
rect 11713 17629 11747 17663
rect 12173 17629 12207 17663
rect 14335 17629 14369 17663
rect 13507 17595 13541 17629
rect 14470 17623 14504 17657
rect 14565 17626 14599 17660
rect 14749 17629 14783 17663
rect 15025 17629 15059 17663
rect 15393 17629 15427 17663
rect 15668 17629 15702 17663
rect 15761 17629 15795 17663
rect 19625 17629 19659 17663
rect 19717 17629 19751 17663
rect 20545 17629 20579 17663
rect 20634 17629 20668 17663
rect 20729 17626 20763 17660
rect 20913 17629 20947 17663
rect 21833 17629 21867 17663
rect 23121 17629 23155 17663
rect 6254 17561 6288 17595
rect 8033 17561 8067 17595
rect 9198 17561 9232 17595
rect 12633 17561 12667 17595
rect 13277 17561 13311 17595
rect 15945 17561 15979 17595
rect 17724 17561 17758 17595
rect 18613 17561 18647 17595
rect 18797 17561 18831 17595
rect 22017 17561 22051 17595
rect 22477 17561 22511 17595
rect 22937 17561 22971 17595
rect 23765 17561 23799 17595
rect 23949 17561 23983 17595
rect 7389 17493 7423 17527
rect 11897 17493 11931 17527
rect 12833 17493 12867 17527
rect 14105 17493 14139 17527
rect 16221 17493 16255 17527
rect 16589 17493 16623 17527
rect 19257 17493 19291 17527
rect 20269 17493 20303 17527
rect 21649 17493 21683 17527
rect 23581 17493 23615 17527
rect 24501 17493 24535 17527
rect 6009 17289 6043 17323
rect 7021 17289 7055 17323
rect 8677 17289 8711 17323
rect 9873 17289 9907 17323
rect 14749 17289 14783 17323
rect 17509 17289 17543 17323
rect 18705 17289 18739 17323
rect 21005 17289 21039 17323
rect 25329 17289 25363 17323
rect 28181 17289 28215 17323
rect 7389 17221 7423 17255
rect 9781 17221 9815 17255
rect 11774 17221 11808 17255
rect 13185 17221 13219 17255
rect 13369 17221 13403 17255
rect 14933 17221 14967 17255
rect 15117 17221 15151 17255
rect 16957 17221 16991 17255
rect 19892 17221 19926 17255
rect 5825 17153 5859 17187
rect 6377 17153 6411 17187
rect 6561 17153 6595 17187
rect 8493 17153 8527 17187
rect 8953 17153 8987 17187
rect 9137 17153 9171 17187
rect 10701 17153 10735 17187
rect 14105 17153 14139 17187
rect 14197 17153 14231 17187
rect 14289 17153 14323 17187
rect 14473 17153 14507 17187
rect 15393 17153 15427 17187
rect 17601 17153 17635 17187
rect 18245 17153 18279 17187
rect 18521 17153 18555 17187
rect 19625 17153 19659 17187
rect 21465 17153 21499 17187
rect 22017 17153 22051 17187
rect 22201 17153 22235 17187
rect 23213 17153 23247 17187
rect 24205 17153 24239 17187
rect 27813 17153 27847 17187
rect 28365 17153 28399 17187
rect 6745 17085 6779 17119
rect 7481 17085 7515 17119
rect 7665 17085 7699 17119
rect 9321 17085 9355 17119
rect 10793 17085 10827 17119
rect 10977 17085 11011 17119
rect 11529 17085 11563 17119
rect 15669 17085 15703 17119
rect 17325 17085 17359 17119
rect 23489 17085 23523 17119
rect 23949 17085 23983 17119
rect 1409 17017 1443 17051
rect 10333 16949 10367 16983
rect 12909 16949 12943 16983
rect 13829 16949 13863 16983
rect 17969 16949 18003 16983
rect 18337 16949 18371 16983
rect 19073 16949 19107 16983
rect 21281 16949 21315 16983
rect 21833 16949 21867 16983
rect 7205 16745 7239 16779
rect 10793 16745 10827 16779
rect 11161 16745 11195 16779
rect 12173 16745 12207 16779
rect 16865 16745 16899 16779
rect 17233 16745 17267 16779
rect 19533 16745 19567 16779
rect 20361 16745 20395 16779
rect 23857 16745 23891 16779
rect 25053 16745 25087 16779
rect 14105 16677 14139 16711
rect 14933 16677 14967 16711
rect 16221 16677 16255 16711
rect 22661 16677 22695 16711
rect 8585 16609 8619 16643
rect 9689 16609 9723 16643
rect 9873 16609 9907 16643
rect 12541 16609 12575 16643
rect 14565 16609 14599 16643
rect 15761 16609 15795 16643
rect 16957 16609 16991 16643
rect 18153 16609 18187 16643
rect 24777 16609 24811 16643
rect 28365 16609 28399 16643
rect 1685 16541 1719 16575
rect 10517 16541 10551 16575
rect 10609 16541 10643 16575
rect 11713 16541 11747 16575
rect 12725 16541 12759 16575
rect 13001 16541 13035 16575
rect 13277 16541 13311 16575
rect 13369 16541 13403 16575
rect 13553 16541 13587 16575
rect 14289 16541 14323 16575
rect 14381 16541 14415 16575
rect 14657 16541 14691 16575
rect 15117 16541 15151 16575
rect 15393 16541 15427 16575
rect 15669 16541 15703 16575
rect 15945 16541 15979 16575
rect 16037 16541 16071 16575
rect 17049 16541 17083 16575
rect 18061 16541 18095 16575
rect 18613 16541 18647 16575
rect 19257 16541 19291 16575
rect 19533 16541 19567 16575
rect 20545 16541 20579 16575
rect 21741 16541 21775 16575
rect 21925 16541 21959 16575
rect 22017 16541 22051 16575
rect 22109 16541 22143 16575
rect 23213 16541 23247 16575
rect 23397 16541 23431 16575
rect 23489 16541 23523 16575
rect 23581 16541 23615 16575
rect 8318 16473 8352 16507
rect 11253 16473 11287 16507
rect 11897 16473 11931 16507
rect 15301 16473 15335 16507
rect 16773 16473 16807 16507
rect 20729 16473 20763 16507
rect 21189 16473 21223 16507
rect 21373 16473 21407 16507
rect 22845 16473 22879 16507
rect 24409 16473 24443 16507
rect 24593 16473 24627 16507
rect 1501 16405 1535 16439
rect 9229 16405 9263 16439
rect 9597 16405 9631 16439
rect 12909 16405 12943 16439
rect 13737 16405 13771 16439
rect 17601 16405 17635 16439
rect 17969 16405 18003 16439
rect 18797 16405 18831 16439
rect 19809 16405 19843 16439
rect 21005 16405 21039 16439
rect 22385 16405 22419 16439
rect 7665 16201 7699 16235
rect 12843 16201 12877 16235
rect 16773 16201 16807 16235
rect 20269 16201 20303 16235
rect 25329 16201 25363 16235
rect 12633 16133 12667 16167
rect 13277 16133 13311 16167
rect 17049 16133 17083 16167
rect 19441 16133 19475 16167
rect 23673 16133 23707 16167
rect 24194 16133 24228 16167
rect 13507 16099 13541 16133
rect 5825 16065 5859 16099
rect 6009 16065 6043 16099
rect 6653 16065 6687 16099
rect 6823 16055 6857 16089
rect 8769 16065 8803 16099
rect 8861 16065 8895 16099
rect 9588 16065 9622 16099
rect 11161 16065 11195 16099
rect 11897 16065 11931 16099
rect 14013 16065 14047 16099
rect 14289 16065 14323 16099
rect 14381 16065 14415 16099
rect 14565 16065 14599 16099
rect 14841 16065 14875 16099
rect 15117 16065 15151 16099
rect 15209 16065 15243 16099
rect 16037 16065 16071 16099
rect 16313 16065 16347 16099
rect 17233 16065 17267 16099
rect 17417 16065 17451 16099
rect 17601 16065 17635 16099
rect 17877 16065 17911 16099
rect 18337 16065 18371 16099
rect 18889 16065 18923 16099
rect 19809 16065 19843 16099
rect 19993 16065 20027 16099
rect 20085 16065 20119 16099
rect 20913 16065 20947 16099
rect 21005 16065 21039 16099
rect 21097 16065 21131 16099
rect 21281 16065 21315 16099
rect 21833 16065 21867 16099
rect 22017 16065 22051 16099
rect 22109 16065 22143 16099
rect 22201 16065 22235 16099
rect 23029 16065 23063 16099
rect 23208 16065 23242 16099
rect 23308 16065 23342 16099
rect 23397 16065 23431 16099
rect 25605 16065 25639 16099
rect 7757 15997 7791 16031
rect 7849 15997 7883 16031
rect 9321 15997 9355 16031
rect 11989 15997 12023 16031
rect 12081 15997 12115 16031
rect 14105 15997 14139 16031
rect 14933 15997 14967 16031
rect 16129 15997 16163 16031
rect 18981 15997 19015 16031
rect 23949 15997 23983 16031
rect 7297 15929 7331 15963
rect 13001 15929 13035 15963
rect 13645 15929 13679 15963
rect 15393 15929 15427 15963
rect 15853 15929 15887 15963
rect 19441 15929 19475 15963
rect 5641 15861 5675 15895
rect 7021 15861 7055 15895
rect 9045 15861 9079 15895
rect 10701 15861 10735 15895
rect 10977 15861 11011 15895
rect 11529 15861 11563 15895
rect 12817 15861 12851 15895
rect 13461 15861 13495 15895
rect 16313 15861 16347 15895
rect 18705 15861 18739 15895
rect 19809 15861 19843 15895
rect 20637 15861 20671 15895
rect 22477 15861 22511 15895
rect 7297 15657 7331 15691
rect 8309 15657 8343 15691
rect 9689 15657 9723 15691
rect 11713 15657 11747 15691
rect 13553 15657 13587 15691
rect 13737 15657 13771 15691
rect 22109 15657 22143 15691
rect 24041 15657 24075 15691
rect 7021 15589 7055 15623
rect 20545 15589 20579 15623
rect 21097 15589 21131 15623
rect 7849 15521 7883 15555
rect 11069 15521 11103 15555
rect 13093 15521 13127 15555
rect 14105 15521 14139 15555
rect 17877 15521 17911 15555
rect 19533 15521 19567 15555
rect 20361 15521 20395 15555
rect 21465 15521 21499 15555
rect 24409 15521 24443 15555
rect 5181 15453 5215 15487
rect 5641 15453 5675 15487
rect 7665 15453 7699 15487
rect 7757 15453 7791 15487
rect 8493 15453 8527 15487
rect 9505 15453 9539 15487
rect 11253 15453 11287 15487
rect 15853 15453 15887 15487
rect 18153 15453 18187 15487
rect 19257 15453 19291 15487
rect 21281 15453 21315 15487
rect 22385 15453 22419 15487
rect 22569 15453 22603 15487
rect 23035 15453 23069 15487
rect 13599 15419 13633 15453
rect 23208 15447 23242 15481
rect 23305 15453 23339 15487
rect 23417 15453 23451 15487
rect 28365 15453 28399 15487
rect 5886 15385 5920 15419
rect 11437 15385 11471 15419
rect 12826 15385 12860 15419
rect 13369 15385 13403 15419
rect 14372 15385 14406 15419
rect 20821 15385 20855 15419
rect 21741 15385 21775 15419
rect 21925 15385 21959 15419
rect 23673 15385 23707 15419
rect 24654 15385 24688 15419
rect 5365 15317 5399 15351
rect 15485 15317 15519 15351
rect 17141 15317 17175 15351
rect 22753 15317 22787 15351
rect 25789 15317 25823 15351
rect 10885 15113 10919 15147
rect 12541 15113 12575 15147
rect 15025 15113 15059 15147
rect 16313 15113 16347 15147
rect 17785 15113 17819 15147
rect 19441 15113 19475 15147
rect 19901 15113 19935 15147
rect 21281 15113 21315 15147
rect 22017 15113 22051 15147
rect 25145 15113 25179 15147
rect 9750 15045 9784 15079
rect 12817 15045 12851 15079
rect 20053 15045 20087 15079
rect 20269 15045 20303 15079
rect 23581 15045 23615 15079
rect 24869 15045 24903 15079
rect 7849 14977 7883 15011
rect 8116 14977 8150 15011
rect 9505 14977 9539 15011
rect 11805 14977 11839 15011
rect 12357 14977 12391 15011
rect 13553 14977 13587 15011
rect 13737 14977 13771 15011
rect 15301 14977 15335 15011
rect 15393 14977 15427 15011
rect 15485 14977 15519 15011
rect 15669 14977 15703 15011
rect 16129 14977 16163 15011
rect 16313 14977 16347 15011
rect 16773 14977 16807 15011
rect 16957 14977 16991 15011
rect 17233 14977 17267 15011
rect 17417 14977 17451 15011
rect 18245 14977 18279 15011
rect 19073 14977 19107 15011
rect 20729 14977 20763 15011
rect 20913 14977 20947 15011
rect 21373 14977 21407 15011
rect 21833 14977 21867 15011
rect 22569 14977 22603 15011
rect 23765 14977 23799 15011
rect 16681 14909 16715 14943
rect 20545 14909 20579 14943
rect 22293 14909 22327 14943
rect 23397 14909 23431 14943
rect 14381 14841 14415 14875
rect 19625 14841 19659 14875
rect 24409 14841 24443 14875
rect 9229 14773 9263 14807
rect 11897 14773 11931 14807
rect 13277 14773 13311 14807
rect 13645 14773 13679 14807
rect 14749 14773 14783 14807
rect 17969 14773 18003 14807
rect 18521 14773 18555 14807
rect 19441 14773 19475 14807
rect 20085 14773 20119 14807
rect 24041 14773 24075 14807
rect 13093 14569 13127 14603
rect 15117 14569 15151 14603
rect 16037 14569 16071 14603
rect 19441 14569 19475 14603
rect 19625 14569 19659 14603
rect 21373 14569 21407 14603
rect 22569 14569 22603 14603
rect 23029 14569 23063 14603
rect 7941 14501 7975 14535
rect 13645 14501 13679 14535
rect 16865 14501 16899 14535
rect 18797 14501 18831 14535
rect 14105 14433 14139 14467
rect 15945 14433 15979 14467
rect 16129 14433 16163 14467
rect 19349 14433 19383 14467
rect 19993 14433 20027 14467
rect 22201 14433 22235 14467
rect 6561 14365 6595 14399
rect 9137 14365 9171 14399
rect 11345 14365 11379 14399
rect 13277 14365 13311 14399
rect 13553 14365 13587 14399
rect 14381 14365 14415 14399
rect 14473 14365 14507 14399
rect 14565 14365 14599 14399
rect 14749 14365 14783 14399
rect 15301 14365 15335 14399
rect 16313 14365 16347 14399
rect 16773 14365 16807 14399
rect 16957 14365 16991 14399
rect 17049 14365 17083 14399
rect 17693 14365 17727 14399
rect 18061 14365 18095 14399
rect 18178 14365 18212 14399
rect 18613 14365 18647 14399
rect 19257 14365 19291 14399
rect 20177 14365 20211 14399
rect 20637 14365 20671 14399
rect 21189 14365 21223 14399
rect 21833 14365 21867 14399
rect 22017 14365 22051 14399
rect 22477 14365 22511 14399
rect 22661 14365 22695 14399
rect 22937 14365 22971 14399
rect 23121 14365 23155 14399
rect 23581 14365 23615 14399
rect 23857 14365 23891 14399
rect 25789 14365 25823 14399
rect 26065 14365 26099 14399
rect 6828 14297 6862 14331
rect 11612 14297 11646 14331
rect 15485 14297 15519 14331
rect 17969 14297 18003 14331
rect 20821 14297 20855 14331
rect 25522 14297 25556 14331
rect 26310 14297 26344 14331
rect 9045 14229 9079 14263
rect 9505 14229 9539 14263
rect 12725 14229 12759 14263
rect 16221 14229 16255 14263
rect 18337 14229 18371 14263
rect 20361 14229 20395 14263
rect 23397 14229 23431 14263
rect 24041 14229 24075 14263
rect 24409 14229 24443 14263
rect 27445 14229 27479 14263
rect 6929 14025 6963 14059
rect 8217 14025 8251 14059
rect 13185 14025 13219 14059
rect 16221 14025 16255 14059
rect 18613 14025 18647 14059
rect 25789 14025 25823 14059
rect 26065 14025 26099 14059
rect 26433 14025 26467 14059
rect 6653 13957 6687 13991
rect 9137 13957 9171 13991
rect 12449 13957 12483 13991
rect 13461 13957 13495 13991
rect 14626 13957 14660 13991
rect 18153 13957 18187 13991
rect 19533 13957 19567 13991
rect 20085 13957 20119 13991
rect 20545 13957 20579 13991
rect 22968 13957 23002 13991
rect 4896 13889 4930 13923
rect 7113 13889 7147 13923
rect 7573 13889 7607 13923
rect 8493 13889 8527 13923
rect 8585 13889 8619 13923
rect 8953 13889 8987 13923
rect 9229 13889 9263 13923
rect 9761 13889 9795 13923
rect 11713 13889 11747 13923
rect 12173 13889 12207 13923
rect 12266 13889 12300 13923
rect 12541 13889 12575 13923
rect 12679 13889 12713 13923
rect 13737 13889 13771 13923
rect 13829 13889 13863 13923
rect 13921 13889 13955 13923
rect 14105 13889 14139 13923
rect 16129 13889 16163 13923
rect 16957 13889 16991 13923
rect 17785 13889 17819 13923
rect 18429 13889 18463 13923
rect 18613 13889 18647 13923
rect 18981 13889 19015 13923
rect 20637 13889 20671 13923
rect 20913 13889 20947 13923
rect 21097 13889 21131 13923
rect 24041 13889 24075 13923
rect 24133 13889 24167 13923
rect 24961 13889 24995 13923
rect 25605 13889 25639 13923
rect 27813 13889 27847 13923
rect 28273 13889 28307 13923
rect 1409 13821 1443 13855
rect 4629 13821 4663 13855
rect 7481 13821 7515 13855
rect 9505 13821 9539 13855
rect 14381 13821 14415 13855
rect 16681 13821 16715 13855
rect 23213 13821 23247 13855
rect 24225 13821 24259 13855
rect 24777 13821 24811 13855
rect 28089 13821 28123 13855
rect 6009 13753 6043 13787
rect 11805 13753 11839 13787
rect 17877 13753 17911 13787
rect 8217 13685 8251 13719
rect 8309 13685 8343 13719
rect 8401 13685 8435 13719
rect 9045 13685 9079 13719
rect 10885 13685 10919 13719
rect 12817 13685 12851 13719
rect 15761 13685 15795 13719
rect 17969 13685 18003 13719
rect 18153 13685 18187 13719
rect 18981 13685 19015 13719
rect 19993 13685 20027 13719
rect 21833 13685 21867 13719
rect 23673 13685 23707 13719
rect 25145 13685 25179 13719
rect 6285 13481 6319 13515
rect 6561 13481 6595 13515
rect 7205 13481 7239 13515
rect 7389 13481 7423 13515
rect 9597 13481 9631 13515
rect 10057 13481 10091 13515
rect 11345 13481 11379 13515
rect 14197 13481 14231 13515
rect 14933 13481 14967 13515
rect 15485 13481 15519 13515
rect 16589 13481 16623 13515
rect 18705 13481 18739 13515
rect 22201 13481 22235 13515
rect 23857 13481 23891 13515
rect 25237 13481 25271 13515
rect 6469 13413 6503 13447
rect 14565 13413 14599 13447
rect 16221 13413 16255 13447
rect 6653 13345 6687 13379
rect 8033 13345 8067 13379
rect 10885 13345 10919 13379
rect 13461 13345 13495 13379
rect 16497 13345 16531 13379
rect 21005 13345 21039 13379
rect 22753 13345 22787 13379
rect 24593 13345 24627 13379
rect 6745 13277 6779 13311
rect 6929 13277 6963 13311
rect 8953 13277 8987 13311
rect 9137 13277 9171 13311
rect 9229 13277 9263 13311
rect 9321 13277 9355 13311
rect 10977 13277 11011 13311
rect 12449 13277 12483 13311
rect 12597 13277 12631 13311
rect 12725 13277 12759 13311
rect 12955 13277 12989 13311
rect 13369 13277 13403 13311
rect 14105 13277 14139 13311
rect 14289 13277 14323 13311
rect 15761 13277 15795 13311
rect 16405 13277 16439 13311
rect 16681 13277 16715 13311
rect 17233 13277 17267 13311
rect 17417 13277 17451 13311
rect 17509 13277 17543 13311
rect 17601 13277 17635 13311
rect 18245 13277 18279 13311
rect 18613 13277 18647 13311
rect 18889 13277 18923 13311
rect 19257 13277 19291 13311
rect 19533 13277 19567 13311
rect 20545 13277 20579 13311
rect 21189 13277 21223 13311
rect 21557 13277 21591 13311
rect 22569 13277 22603 13311
rect 23489 13277 23523 13311
rect 23673 13277 23707 13311
rect 25513 13277 25547 13311
rect 7573 13209 7607 13243
rect 8309 13209 8343 13243
rect 8585 13209 8619 13243
rect 10241 13209 10275 13243
rect 12817 13209 12851 13243
rect 20361 13209 20395 13243
rect 25758 13209 25792 13243
rect 7373 13141 7407 13175
rect 8217 13141 8251 13175
rect 8401 13141 8435 13175
rect 9873 13141 9907 13175
rect 10041 13141 10075 13175
rect 13093 13141 13127 13175
rect 15945 13141 15979 13175
rect 17877 13141 17911 13175
rect 18429 13141 18463 13175
rect 20729 13141 20763 13175
rect 21741 13141 21775 13175
rect 22661 13141 22695 13175
rect 24777 13141 24811 13175
rect 24869 13141 24903 13175
rect 26893 13141 26927 13175
rect 7005 12937 7039 12971
rect 7481 12937 7515 12971
rect 7941 12937 7975 12971
rect 13185 12937 13219 12971
rect 15669 12937 15703 12971
rect 17141 12937 17175 12971
rect 18337 12937 18371 12971
rect 19441 12937 19475 12971
rect 24041 12937 24075 12971
rect 25605 12937 25639 12971
rect 7205 12869 7239 12903
rect 8921 12869 8955 12903
rect 9137 12869 9171 12903
rect 13737 12869 13771 12903
rect 14381 12869 14415 12903
rect 16773 12869 16807 12903
rect 24777 12869 24811 12903
rect 26341 12869 26375 12903
rect 4445 12801 4479 12835
rect 4712 12801 4746 12835
rect 7481 12801 7515 12835
rect 7665 12801 7699 12835
rect 8125 12801 8159 12835
rect 8309 12801 8343 12835
rect 11713 12801 11747 12835
rect 12817 12801 12851 12835
rect 13277 12801 13311 12835
rect 14565 12801 14599 12835
rect 14841 12801 14875 12835
rect 15025 12801 15059 12835
rect 16037 12801 16071 12835
rect 16129 12801 16163 12835
rect 16957 12801 16991 12835
rect 17417 12801 17451 12835
rect 17601 12801 17635 12835
rect 18245 12801 18279 12835
rect 18429 12801 18463 12835
rect 19165 12801 19199 12835
rect 19625 12801 19659 12835
rect 19809 12801 19843 12835
rect 20352 12801 20386 12835
rect 21925 12801 21959 12835
rect 22652 12801 22686 12835
rect 25421 12801 25455 12835
rect 26065 12801 26099 12835
rect 8217 12733 8251 12767
rect 8401 12733 8435 12767
rect 9689 12733 9723 12767
rect 9965 12733 9999 12767
rect 11621 12733 11655 12767
rect 12081 12733 12115 12767
rect 13921 12733 13955 12767
rect 15209 12733 15243 12767
rect 20085 12733 20119 12767
rect 22385 12733 22419 12767
rect 24869 12733 24903 12767
rect 24961 12733 24995 12767
rect 8769 12665 8803 12699
rect 22109 12665 22143 12699
rect 5825 12597 5859 12631
rect 6837 12597 6871 12631
rect 7021 12597 7055 12631
rect 8953 12597 8987 12631
rect 10977 12597 11011 12631
rect 14197 12597 14231 12631
rect 16313 12597 16347 12631
rect 17785 12597 17819 12631
rect 18705 12597 18739 12631
rect 18889 12597 18923 12631
rect 21465 12597 21499 12631
rect 23765 12597 23799 12631
rect 24409 12597 24443 12631
rect 25881 12597 25915 12631
rect 28365 12597 28399 12631
rect 5549 12393 5583 12427
rect 6745 12393 6779 12427
rect 8585 12393 8619 12427
rect 9137 12393 9171 12427
rect 9965 12393 9999 12427
rect 10609 12393 10643 12427
rect 12357 12393 12391 12427
rect 20453 12393 20487 12427
rect 23489 12393 23523 12427
rect 24777 12393 24811 12427
rect 10333 12257 10367 12291
rect 11989 12257 12023 12291
rect 21097 12257 21131 12291
rect 22753 12257 22787 12291
rect 24409 12257 24443 12291
rect 5825 12189 5859 12223
rect 5917 12189 5951 12223
rect 6009 12189 6043 12223
rect 6193 12189 6227 12223
rect 7941 12189 7975 12223
rect 8309 12189 8343 12223
rect 8585 12189 8619 12223
rect 10149 12189 10183 12223
rect 13737 12189 13771 12223
rect 14473 12189 14507 12223
rect 14565 12189 14599 12223
rect 14657 12189 14691 12223
rect 14841 12189 14875 12223
rect 15393 12189 15427 12223
rect 15485 12189 15519 12223
rect 15577 12189 15611 12223
rect 15761 12189 15795 12223
rect 16037 12189 16071 12223
rect 16129 12189 16163 12223
rect 16313 12189 16347 12223
rect 16405 12189 16439 12223
rect 17141 12189 17175 12223
rect 17325 12189 17359 12223
rect 17417 12189 17451 12223
rect 17509 12189 17543 12223
rect 19717 12189 19751 12223
rect 20821 12189 20855 12223
rect 21649 12189 21683 12223
rect 21741 12189 21775 12223
rect 23305 12189 23339 12223
rect 24041 12189 24075 12223
rect 24593 12189 24627 12223
rect 25421 12189 25455 12223
rect 6561 12121 6595 12155
rect 6761 12121 6795 12155
rect 7481 12121 7515 12155
rect 8493 12121 8527 12155
rect 9105 12121 9139 12155
rect 9321 12121 9355 12155
rect 11722 12121 11756 12155
rect 13492 12121 13526 12155
rect 15117 12121 15151 12155
rect 19901 12121 19935 12155
rect 22569 12121 22603 12155
rect 25053 12121 25087 12155
rect 25688 12121 25722 12155
rect 6929 12053 6963 12087
rect 7573 12053 7607 12087
rect 8953 12053 8987 12087
rect 14197 12053 14231 12087
rect 16589 12053 16623 12087
rect 17785 12053 17819 12087
rect 18245 12053 18279 12087
rect 18613 12053 18647 12087
rect 19349 12053 19383 12087
rect 20913 12053 20947 12087
rect 21925 12053 21959 12087
rect 22201 12053 22235 12087
rect 22661 12053 22695 12087
rect 23857 12053 23891 12087
rect 26801 12053 26835 12087
rect 10885 11849 10919 11883
rect 13001 11849 13035 11883
rect 15853 11849 15887 11883
rect 18337 11849 18371 11883
rect 20453 11849 20487 11883
rect 21097 11849 21131 11883
rect 23029 11849 23063 11883
rect 24501 11849 24535 11883
rect 25973 11849 26007 11883
rect 5273 11781 5307 11815
rect 5825 11781 5859 11815
rect 6929 11781 6963 11815
rect 14350 11781 14384 11815
rect 17794 11781 17828 11815
rect 20545 11781 20579 11815
rect 23581 11781 23615 11815
rect 23765 11781 23799 11815
rect 28089 11781 28123 11815
rect 5365 11713 5399 11747
rect 5641 11713 5675 11747
rect 5917 11713 5951 11747
rect 6745 11713 6779 11747
rect 6837 11713 6871 11747
rect 7113 11713 7147 11747
rect 7205 11713 7239 11747
rect 7757 11713 7791 11747
rect 9321 11713 9355 11747
rect 9781 11713 9815 11747
rect 9965 11713 9999 11747
rect 10241 11713 10275 11747
rect 10425 11713 10459 11747
rect 10520 11716 10554 11750
rect 10609 11713 10643 11747
rect 12081 11713 12115 11747
rect 12541 11713 12575 11747
rect 12725 11713 12759 11747
rect 14105 11713 14139 11747
rect 15945 11713 15979 11747
rect 18797 11713 18831 11747
rect 19533 11713 19567 11747
rect 21281 11713 21315 11747
rect 22109 11713 22143 11747
rect 22753 11713 22787 11747
rect 23213 11713 23247 11747
rect 24593 11713 24627 11747
rect 27813 11713 27847 11747
rect 28273 11713 28307 11747
rect 8033 11645 8067 11679
rect 9229 11645 9263 11679
rect 18061 11645 18095 11679
rect 20637 11645 20671 11679
rect 22293 11645 22327 11679
rect 24777 11645 24811 11679
rect 26065 11645 26099 11679
rect 26157 11645 26191 11679
rect 6561 11577 6595 11611
rect 11621 11577 11655 11611
rect 16681 11577 16715 11611
rect 5641 11509 5675 11543
rect 8953 11509 8987 11543
rect 9781 11509 9815 11543
rect 12173 11509 12207 11543
rect 12633 11509 12667 11543
rect 13829 11509 13863 11543
rect 15485 11509 15519 11543
rect 18981 11509 19015 11543
rect 19349 11509 19383 11543
rect 20085 11509 20119 11543
rect 22569 11509 22603 11543
rect 24133 11509 24167 11543
rect 25605 11509 25639 11543
rect 4537 11305 4571 11339
rect 6837 11305 6871 11339
rect 7297 11305 7331 11339
rect 8585 11305 8619 11339
rect 9643 11305 9677 11339
rect 9873 11305 9907 11339
rect 12541 11305 12575 11339
rect 12633 11305 12667 11339
rect 15117 11305 15151 11339
rect 15761 11305 15795 11339
rect 17049 11305 17083 11339
rect 19349 11305 19383 11339
rect 21005 11305 21039 11339
rect 24409 11305 24443 11339
rect 25513 11305 25547 11339
rect 7665 11237 7699 11271
rect 12449 11237 12483 11271
rect 13645 11237 13679 11271
rect 14381 11237 14415 11271
rect 14749 11237 14783 11271
rect 16497 11237 16531 11271
rect 23857 11237 23891 11271
rect 27169 11237 27203 11271
rect 7021 11169 7055 11203
rect 11805 11169 11839 11203
rect 15025 11169 15059 11203
rect 23305 11169 23339 11203
rect 23397 11169 23431 11203
rect 24869 11169 24903 11203
rect 25053 11169 25087 11203
rect 5917 11101 5951 11135
rect 7113 11101 7147 11135
rect 7573 11101 7607 11135
rect 7757 11101 7791 11135
rect 8125 11101 8159 11135
rect 8217 11101 8251 11135
rect 8401 11101 8435 11135
rect 9137 11101 9171 11135
rect 9505 11101 9539 11135
rect 9781 11101 9815 11135
rect 9965 11101 9999 11135
rect 10609 11101 10643 11135
rect 10793 11101 10827 11135
rect 10885 11101 10919 11135
rect 10977 11101 11011 11135
rect 12357 11101 12391 11135
rect 12817 11101 12851 11135
rect 13093 11101 13127 11135
rect 13277 11101 13311 11135
rect 13461 11101 13495 11135
rect 14933 11101 14967 11135
rect 16681 11101 16715 11135
rect 18797 11101 18831 11135
rect 19625 11101 19659 11135
rect 21373 11101 21407 11135
rect 25145 11101 25179 11135
rect 25789 11101 25823 11135
rect 5650 11033 5684 11067
rect 6837 11033 6871 11067
rect 8953 11033 8987 11067
rect 11621 11033 11655 11067
rect 13369 11033 13403 11067
rect 14197 11033 14231 11067
rect 15209 11033 15243 11067
rect 16129 11033 16163 11067
rect 18530 11033 18564 11067
rect 19870 11033 19904 11067
rect 21640 11033 21674 11067
rect 23489 11033 23523 11067
rect 26056 11033 26090 11067
rect 11253 10965 11287 10999
rect 12081 10965 12115 10999
rect 17417 10965 17451 10999
rect 22753 10965 22787 10999
rect 7849 10761 7883 10795
rect 8861 10761 8895 10795
rect 10885 10761 10919 10795
rect 16957 10761 16991 10795
rect 17509 10761 17543 10795
rect 19257 10761 19291 10795
rect 20729 10761 20763 10795
rect 25789 10761 25823 10795
rect 26433 10761 26467 10795
rect 9382 10693 9416 10727
rect 11774 10693 11808 10727
rect 14473 10693 14507 10727
rect 14657 10693 14691 10727
rect 15025 10693 15059 10727
rect 17049 10693 17083 10727
rect 18622 10693 18656 10727
rect 19349 10693 19383 10727
rect 21373 10693 21407 10727
rect 22477 10693 22511 10727
rect 23756 10693 23790 10727
rect 5641 10625 5675 10659
rect 6653 10625 6687 10659
rect 6837 10625 6871 10659
rect 7113 10625 7147 10659
rect 7389 10625 7423 10659
rect 7757 10625 7791 10659
rect 8677 10625 8711 10659
rect 9137 10625 9171 10659
rect 10793 10625 10827 10659
rect 10977 10625 11011 10659
rect 11529 10625 11563 10659
rect 13461 10625 13495 10659
rect 15301 10625 15335 10659
rect 18889 10625 18923 10659
rect 19901 10625 19935 10659
rect 20085 10625 20119 10659
rect 20361 10625 20395 10659
rect 20545 10625 20579 10659
rect 21005 10625 21039 10659
rect 22385 10625 22419 10659
rect 23213 10625 23247 10659
rect 23489 10625 23523 10659
rect 26617 10625 26651 10659
rect 28089 10625 28123 10659
rect 13185 10557 13219 10591
rect 15209 10557 15243 10591
rect 22569 10557 22603 10591
rect 25513 10557 25547 10591
rect 25697 10557 25731 10591
rect 7389 10489 7423 10523
rect 12909 10489 12943 10523
rect 24869 10489 24903 10523
rect 1409 10421 1443 10455
rect 5457 10421 5491 10455
rect 6837 10421 6871 10455
rect 8309 10421 8343 10455
rect 10517 10421 10551 10455
rect 14289 10421 14323 10455
rect 15025 10421 15059 10455
rect 15485 10421 15519 10455
rect 19717 10421 19751 10455
rect 22017 10421 22051 10455
rect 23029 10421 23063 10455
rect 26157 10421 26191 10455
rect 28273 10421 28307 10455
rect 7297 10217 7331 10251
rect 8953 10217 8987 10251
rect 13185 10217 13219 10251
rect 13553 10217 13587 10251
rect 22385 10217 22419 10251
rect 25605 10217 25639 10251
rect 6561 10149 6595 10183
rect 15485 10149 15519 10183
rect 17693 10149 17727 10183
rect 7573 10081 7607 10115
rect 9137 10081 9171 10115
rect 9413 10081 9447 10115
rect 11161 10081 11195 10115
rect 11437 10081 11471 10115
rect 14933 10081 14967 10115
rect 15577 10081 15611 10115
rect 19809 10081 19843 10115
rect 21833 10081 21867 10115
rect 21925 10081 21959 10115
rect 24501 10081 24535 10115
rect 5181 10013 5215 10047
rect 6929 10013 6963 10047
rect 7113 10013 7147 10047
rect 7849 10013 7883 10047
rect 9229 10013 9263 10047
rect 9321 10013 9355 10047
rect 12817 10013 12851 10047
rect 13461 10013 13495 10047
rect 13645 10013 13679 10047
rect 14105 10013 14139 10047
rect 14289 10013 14323 10047
rect 14749 10013 14783 10047
rect 15393 10013 15427 10047
rect 15669 10013 15703 10047
rect 16681 10013 16715 10047
rect 17049 10013 17083 10047
rect 17417 10013 17451 10047
rect 18337 10013 18371 10047
rect 18705 10013 18739 10047
rect 19349 10013 19383 10047
rect 22661 10013 22695 10047
rect 24777 10013 24811 10047
rect 26985 10013 27019 10047
rect 27445 10013 27479 10047
rect 5448 9945 5482 9979
rect 12449 9945 12483 9979
rect 13001 9945 13035 9979
rect 14565 9945 14599 9979
rect 18153 9945 18187 9979
rect 20054 9945 20088 9979
rect 22928 9945 22962 9979
rect 26740 9945 26774 9979
rect 12357 9877 12391 9911
rect 14289 9877 14323 9911
rect 15209 9877 15243 9911
rect 16037 9877 16071 9911
rect 17877 9877 17911 9911
rect 19533 9877 19567 9911
rect 21189 9877 21223 9911
rect 22017 9877 22051 9911
rect 24041 9877 24075 9911
rect 24685 9877 24719 9911
rect 25145 9877 25179 9911
rect 27261 9877 27295 9911
rect 8519 9673 8553 9707
rect 14749 9673 14783 9707
rect 16773 9673 16807 9707
rect 19901 9673 19935 9707
rect 21833 9673 21867 9707
rect 24041 9673 24075 9707
rect 24685 9673 24719 9707
rect 25145 9673 25179 9707
rect 25973 9673 26007 9707
rect 26433 9673 26467 9707
rect 7941 9605 7975 9639
rect 8309 9605 8343 9639
rect 11897 9605 11931 9639
rect 12265 9605 12299 9639
rect 16221 9605 16255 9639
rect 18306 9605 18340 9639
rect 20361 9605 20395 9639
rect 21465 9605 21499 9639
rect 25053 9605 25087 9639
rect 26065 9605 26099 9639
rect 7205 9537 7239 9571
rect 7481 9537 7515 9571
rect 7849 9537 7883 9571
rect 8033 9537 8067 9571
rect 9045 9537 9079 9571
rect 9229 9537 9263 9571
rect 9772 9537 9806 9571
rect 12081 9537 12115 9571
rect 12541 9537 12575 9571
rect 12725 9537 12759 9571
rect 12817 9537 12851 9571
rect 14013 9537 14047 9571
rect 14473 9537 14507 9571
rect 16129 9537 16163 9571
rect 16313 9537 16347 9571
rect 16681 9537 16715 9571
rect 16865 9537 16899 9571
rect 17325 9537 17359 9571
rect 17417 9537 17451 9571
rect 17601 9537 17635 9571
rect 18061 9537 18095 9571
rect 20269 9537 20303 9571
rect 21281 9537 21315 9571
rect 22946 9537 22980 9571
rect 23213 9537 23247 9571
rect 5825 9469 5859 9503
rect 9505 9469 9539 9503
rect 14105 9469 14139 9503
rect 14565 9469 14599 9503
rect 14749 9469 14783 9503
rect 20545 9469 20579 9503
rect 24133 9469 24167 9503
rect 24317 9469 24351 9503
rect 25237 9469 25271 9503
rect 25789 9469 25823 9503
rect 5549 9401 5583 9435
rect 5365 9333 5399 9367
rect 7021 9333 7055 9367
rect 7389 9333 7423 9367
rect 8493 9333 8527 9367
rect 8677 9333 8711 9367
rect 10885 9333 10919 9367
rect 12541 9333 12575 9367
rect 13645 9333 13679 9367
rect 17601 9333 17635 9367
rect 19441 9333 19475 9367
rect 23673 9333 23707 9367
rect 7389 9129 7423 9163
rect 9965 9129 9999 9163
rect 16681 9129 16715 9163
rect 20453 9129 20487 9163
rect 22109 9129 22143 9163
rect 7849 9061 7883 9095
rect 15301 9061 15335 9095
rect 21741 9061 21775 9095
rect 19717 8993 19751 9027
rect 22385 8993 22419 9027
rect 24961 8993 24995 9027
rect 1869 8925 1903 8959
rect 6009 8925 6043 8959
rect 7665 8925 7699 8959
rect 7987 8925 8021 8959
rect 8125 8925 8159 8959
rect 9965 8925 9999 8959
rect 10241 8925 10275 8959
rect 10701 8925 10735 8959
rect 10885 8925 10919 8959
rect 11009 8925 11043 8959
rect 11161 8925 11195 8959
rect 11253 8925 11287 8959
rect 12173 8925 12207 8959
rect 12440 8925 12474 8959
rect 15025 8925 15059 8959
rect 16865 8925 16899 8959
rect 16957 8925 16991 8959
rect 17141 8925 17175 8959
rect 17233 8925 17267 8959
rect 17509 8925 17543 8959
rect 17776 8925 17810 8959
rect 19349 8925 19383 8959
rect 19901 8925 19935 8959
rect 20361 8925 20395 8959
rect 20545 8925 20579 8959
rect 21649 8925 21683 8959
rect 21833 8925 21867 8959
rect 21925 8925 21959 8959
rect 22661 8925 22695 8959
rect 26065 8925 26099 8959
rect 28365 8925 28399 8959
rect 1685 8857 1719 8891
rect 2145 8857 2179 8891
rect 6276 8857 6310 8891
rect 11621 8857 11655 8891
rect 11805 8857 11839 8891
rect 15117 8857 15151 8891
rect 15301 8857 15335 8891
rect 7665 8789 7699 8823
rect 10149 8789 10183 8823
rect 13553 8789 13587 8823
rect 18889 8789 18923 8823
rect 20085 8789 20119 8823
rect 25145 8789 25179 8823
rect 25237 8789 25271 8823
rect 25605 8789 25639 8823
rect 25881 8789 25915 8823
rect 6837 8585 6871 8619
rect 8033 8585 8067 8619
rect 10425 8585 10459 8619
rect 12725 8585 12759 8619
rect 14105 8585 14139 8619
rect 18061 8585 18095 8619
rect 22477 8585 22511 8619
rect 24869 8585 24903 8619
rect 2053 8517 2087 8551
rect 11805 8517 11839 8551
rect 12173 8517 12207 8551
rect 12357 8517 12391 8551
rect 17693 8517 17727 8551
rect 19165 8517 19199 8551
rect 19349 8517 19383 8551
rect 22661 8517 22695 8551
rect 22845 8517 22879 8551
rect 25504 8517 25538 8551
rect 1685 8449 1719 8483
rect 4896 8449 4930 8483
rect 7113 8449 7147 8483
rect 7849 8449 7883 8483
rect 8125 8449 8159 8483
rect 8401 8449 8435 8483
rect 8668 8449 8702 8483
rect 10057 8449 10091 8483
rect 10195 8449 10229 8483
rect 10517 8449 10551 8483
rect 10793 8449 10827 8483
rect 10885 8449 10919 8483
rect 11529 8449 11563 8483
rect 12081 8449 12115 8483
rect 13093 8449 13127 8483
rect 13277 8449 13311 8483
rect 13461 8449 13495 8483
rect 14289 8449 14323 8483
rect 14473 8449 14507 8483
rect 14565 8449 14599 8483
rect 15200 8449 15234 8483
rect 16865 8449 16899 8483
rect 17325 8449 17359 8483
rect 17509 8449 17543 8483
rect 17969 8449 18003 8483
rect 18153 8449 18187 8483
rect 19984 8449 20018 8483
rect 23756 8449 23790 8483
rect 25237 8449 25271 8483
rect 4629 8381 4663 8415
rect 6837 8381 6871 8415
rect 10333 8381 10367 8415
rect 11805 8381 11839 8415
rect 13001 8381 13035 8415
rect 14381 8381 14415 8415
rect 14933 8381 14967 8415
rect 17049 8381 17083 8415
rect 19717 8381 19751 8415
rect 23489 8381 23523 8415
rect 9781 8313 9815 8347
rect 12357 8313 12391 8347
rect 16313 8313 16347 8347
rect 18705 8313 18739 8347
rect 21097 8313 21131 8347
rect 26617 8313 26651 8347
rect 6009 8245 6043 8279
rect 7021 8245 7055 8279
rect 7665 8245 7699 8279
rect 10793 8245 10827 8279
rect 11161 8245 11195 8279
rect 11621 8245 11655 8279
rect 13185 8245 13219 8279
rect 16681 8245 16715 8279
rect 1409 8041 1443 8075
rect 6377 8041 6411 8075
rect 10701 8041 10735 8075
rect 11529 8041 11563 8075
rect 11989 8041 12023 8075
rect 12449 8041 12483 8075
rect 13277 8041 13311 8075
rect 14289 8041 14323 8075
rect 15117 8041 15151 8075
rect 15485 8041 15519 8075
rect 16221 8041 16255 8075
rect 16497 8041 16531 8075
rect 16957 8041 16991 8075
rect 17969 8041 18003 8075
rect 19257 8041 19291 8075
rect 20085 8041 20119 8075
rect 21189 8041 21223 8075
rect 23765 8041 23799 8075
rect 25329 8041 25363 8075
rect 14105 7973 14139 8007
rect 19717 7973 19751 8007
rect 6101 7905 6135 7939
rect 8125 7905 8159 7939
rect 10517 7905 10551 7939
rect 11713 7905 11747 7939
rect 12541 7905 12575 7939
rect 15577 7905 15611 7939
rect 19349 7905 19383 7939
rect 25881 7905 25915 7939
rect 5825 7837 5859 7871
rect 5917 7837 5951 7871
rect 6561 7837 6595 7871
rect 6883 7837 6917 7871
rect 7021 7837 7055 7871
rect 7573 7837 7607 7871
rect 7757 7837 7791 7871
rect 8033 7837 8067 7871
rect 8217 7837 8251 7871
rect 9597 7837 9631 7871
rect 10057 7837 10091 7871
rect 10425 7837 10459 7871
rect 10701 7837 10735 7871
rect 11529 7837 11563 7871
rect 11805 7837 11839 7871
rect 12265 7837 12299 7871
rect 12357 7837 12391 7871
rect 15301 7837 15335 7871
rect 15853 7837 15887 7871
rect 16497 7837 16531 7871
rect 16589 7837 16623 7871
rect 17049 7837 17083 7871
rect 17141 7837 17175 7871
rect 18705 7837 18739 7871
rect 19533 7837 19567 7871
rect 20269 7837 20303 7871
rect 20453 7837 20487 7871
rect 20545 7837 20579 7871
rect 20821 7837 20855 7871
rect 21281 7837 21315 7871
rect 23029 7837 23063 7871
rect 23581 7837 23615 7871
rect 24409 7837 24443 7871
rect 25789 7837 25823 7871
rect 27905 7837 27939 7871
rect 28365 7837 28399 7871
rect 6653 7769 6687 7803
rect 6745 7769 6779 7803
rect 13369 7769 13403 7803
rect 14273 7769 14307 7803
rect 14473 7769 14507 7803
rect 16865 7769 16899 7803
rect 19257 7769 19291 7803
rect 22762 7769 22796 7803
rect 6101 7701 6135 7735
rect 7665 7701 7699 7735
rect 9965 7701 9999 7735
rect 10885 7701 10919 7735
rect 17325 7701 17359 7735
rect 18337 7701 18371 7735
rect 18797 7701 18831 7735
rect 20913 7701 20947 7735
rect 21005 7701 21039 7735
rect 21281 7701 21315 7735
rect 21649 7701 21683 7735
rect 24501 7701 24535 7735
rect 25697 7701 25731 7735
rect 28181 7701 28215 7735
rect 7481 7497 7515 7531
rect 8769 7497 8803 7531
rect 17417 7497 17451 7531
rect 24133 7497 24167 7531
rect 24593 7497 24627 7531
rect 4896 7429 4930 7463
rect 7849 7429 7883 7463
rect 9321 7429 9355 7463
rect 17233 7429 17267 7463
rect 21005 7429 21039 7463
rect 21833 7429 21867 7463
rect 21925 7429 21959 7463
rect 22661 7429 22695 7463
rect 22877 7429 22911 7463
rect 24501 7429 24535 7463
rect 4629 7361 4663 7395
rect 6377 7361 6411 7395
rect 7665 7361 7699 7395
rect 7757 7361 7791 7395
rect 8033 7361 8067 7395
rect 8677 7361 8711 7395
rect 9781 7361 9815 7395
rect 9965 7361 9999 7395
rect 10333 7361 10367 7395
rect 10609 7361 10643 7395
rect 11805 7361 11839 7395
rect 13369 7361 13403 7395
rect 13645 7361 13679 7395
rect 14749 7361 14783 7395
rect 14841 7361 14875 7395
rect 15025 7361 15059 7395
rect 15117 7361 15151 7395
rect 15853 7361 15887 7395
rect 15945 7361 15979 7395
rect 16129 7361 16163 7395
rect 17509 7361 17543 7395
rect 17785 7361 17819 7395
rect 18041 7361 18075 7395
rect 19625 7361 19659 7395
rect 20821 7361 20855 7395
rect 23397 7361 23431 7395
rect 25329 7361 25363 7395
rect 6653 7293 6687 7327
rect 12265 7293 12299 7327
rect 12541 7293 12575 7327
rect 19901 7293 19935 7327
rect 22201 7293 22235 7327
rect 22293 7293 22327 7327
rect 24685 7293 24719 7327
rect 25513 7293 25547 7327
rect 6009 7225 6043 7259
rect 9137 7225 9171 7259
rect 17233 7225 17267 7259
rect 23581 7225 23615 7259
rect 9873 7157 9907 7191
rect 11897 7157 11931 7191
rect 14565 7157 14599 7191
rect 16129 7157 16163 7191
rect 19165 7157 19199 7191
rect 22109 7157 22143 7191
rect 22845 7157 22879 7191
rect 23029 7157 23063 7191
rect 25145 7157 25179 7191
rect 6929 6953 6963 6987
rect 7297 6953 7331 6987
rect 10333 6953 10367 6987
rect 15485 6953 15519 6987
rect 17601 6953 17635 6987
rect 18429 6953 18463 6987
rect 20545 6953 20579 6987
rect 24041 6953 24075 6987
rect 12173 6885 12207 6919
rect 12265 6885 12299 6919
rect 17969 6885 18003 6919
rect 20085 6885 20119 6919
rect 24961 6885 24995 6919
rect 8953 6817 8987 6851
rect 17693 6817 17727 6851
rect 19349 6817 19383 6851
rect 20913 6817 20947 6851
rect 22201 6817 22235 6851
rect 6653 6749 6687 6783
rect 6929 6749 6963 6783
rect 7021 6749 7055 6783
rect 7941 6749 7975 6783
rect 8033 6749 8067 6783
rect 8217 6749 8251 6783
rect 8309 6749 8343 6783
rect 10793 6749 10827 6783
rect 10885 6749 10919 6783
rect 11069 6749 11103 6783
rect 11161 6749 11195 6783
rect 11529 6749 11563 6783
rect 12081 6749 12115 6783
rect 12393 6749 12427 6783
rect 12909 6749 12943 6783
rect 13645 6749 13679 6783
rect 14105 6749 14139 6783
rect 15761 6749 15795 6783
rect 16028 6749 16062 6783
rect 17417 6749 17451 6783
rect 17509 6749 17543 6783
rect 18245 6749 18279 6783
rect 18337 6749 18371 6783
rect 18521 6749 18555 6783
rect 18705 6749 18739 6783
rect 19257 6749 19291 6783
rect 19441 6749 19475 6783
rect 21097 6749 21131 6783
rect 21281 6749 21315 6783
rect 21373 6749 21407 6783
rect 21833 6749 21867 6783
rect 22661 6749 22695 6783
rect 25237 6749 25271 6783
rect 6386 6681 6420 6715
rect 9220 6681 9254 6715
rect 14350 6681 14384 6715
rect 19717 6681 19751 6715
rect 21649 6681 21683 6715
rect 22928 6681 22962 6715
rect 24777 6681 24811 6715
rect 25504 6681 25538 6715
rect 5273 6613 5307 6647
rect 7757 6613 7791 6647
rect 10609 6613 10643 6647
rect 11897 6613 11931 6647
rect 12817 6613 12851 6647
rect 13553 6613 13587 6647
rect 17141 6613 17175 6647
rect 20177 6613 20211 6647
rect 26617 6613 26651 6647
rect 6469 6409 6503 6443
rect 8401 6409 8435 6443
rect 8769 6409 8803 6443
rect 9873 6409 9907 6443
rect 13553 6409 13587 6443
rect 14203 6409 14237 6443
rect 14289 6409 14323 6443
rect 14841 6409 14875 6443
rect 16313 6409 16347 6443
rect 21005 6409 21039 6443
rect 23305 6409 23339 6443
rect 25697 6409 25731 6443
rect 6745 6341 6779 6375
rect 6975 6341 7009 6375
rect 8033 6341 8067 6375
rect 8249 6341 8283 6375
rect 11621 6341 11655 6375
rect 17877 6341 17911 6375
rect 19809 6341 19843 6375
rect 20269 6341 20303 6375
rect 22937 6341 22971 6375
rect 25329 6341 25363 6375
rect 25421 6341 25455 6375
rect 6653 6273 6687 6307
rect 6837 6273 6871 6307
rect 7113 6273 7147 6307
rect 7389 6273 7423 6307
rect 7573 6273 7607 6307
rect 8861 6273 8895 6307
rect 9689 6273 9723 6307
rect 9965 6273 9999 6307
rect 10977 6273 11011 6307
rect 11161 6273 11195 6307
rect 12429 6273 12463 6307
rect 14105 6273 14139 6307
rect 14381 6273 14415 6307
rect 14841 6273 14875 6307
rect 15025 6273 15059 6307
rect 16037 6273 16071 6307
rect 16129 6273 16163 6307
rect 18153 6273 18187 6307
rect 18337 6273 18371 6307
rect 19073 6273 19107 6307
rect 19165 6273 19199 6307
rect 19349 6273 19383 6307
rect 20453 6273 20487 6307
rect 20545 6273 20579 6307
rect 20913 6273 20947 6307
rect 22201 6273 22235 6307
rect 23121 6273 23155 6307
rect 23397 6273 23431 6307
rect 23857 6273 23891 6307
rect 24685 6273 24719 6307
rect 25145 6273 25179 6307
rect 25513 6273 25547 6307
rect 12173 6205 12207 6239
rect 16313 6205 16347 6239
rect 21281 6205 21315 6239
rect 21833 6205 21867 6239
rect 22109 6205 22143 6239
rect 23029 6205 23063 6239
rect 7389 6137 7423 6171
rect 9689 6137 9723 6171
rect 11805 6137 11839 6171
rect 18889 6137 18923 6171
rect 19993 6137 20027 6171
rect 21189 6137 21223 6171
rect 24869 6137 24903 6171
rect 8217 6069 8251 6103
rect 10977 6069 11011 6103
rect 18245 6069 18279 6103
rect 19073 6069 19107 6103
rect 20361 6069 20395 6103
rect 21097 6069 21131 6103
rect 24041 6069 24075 6103
rect 8493 5865 8527 5899
rect 12173 5865 12207 5899
rect 13277 5865 13311 5899
rect 14381 5865 14415 5899
rect 14565 5865 14599 5899
rect 18337 5865 18371 5899
rect 19441 5865 19475 5899
rect 21741 5865 21775 5899
rect 22201 5865 22235 5899
rect 22477 5865 22511 5899
rect 23581 5865 23615 5899
rect 9229 5797 9263 5831
rect 14933 5797 14967 5831
rect 16865 5797 16899 5831
rect 21373 5797 21407 5831
rect 22845 5797 22879 5831
rect 23305 5797 23339 5831
rect 8125 5729 8159 5763
rect 9321 5729 9355 5763
rect 13369 5729 13403 5763
rect 18153 5729 18187 5763
rect 19349 5729 19383 5763
rect 19993 5729 20027 5763
rect 24961 5729 24995 5763
rect 1685 5661 1719 5695
rect 7869 5661 7903 5695
rect 9045 5661 9079 5695
rect 9137 5661 9171 5695
rect 9781 5661 9815 5695
rect 9873 5661 9907 5695
rect 10057 5661 10091 5695
rect 10149 5661 10183 5695
rect 10877 5661 10911 5695
rect 10969 5661 11003 5695
rect 11161 5661 11195 5695
rect 11263 5661 11297 5695
rect 11529 5661 11563 5695
rect 11713 5661 11747 5695
rect 11805 5661 11839 5695
rect 11943 5661 11977 5695
rect 13553 5661 13587 5695
rect 16589 5661 16623 5695
rect 16681 5661 16715 5695
rect 17417 5661 17451 5695
rect 17693 5661 17727 5695
rect 18337 5661 18371 5695
rect 19257 5661 19291 5695
rect 20260 5661 20294 5695
rect 21925 5661 21959 5695
rect 22017 5661 22051 5695
rect 22477 5661 22511 5695
rect 22661 5661 22695 5695
rect 23765 5661 23799 5695
rect 24777 5661 24811 5695
rect 28365 5661 28399 5695
rect 12633 5593 12667 5627
rect 13277 5593 13311 5627
rect 14565 5593 14599 5627
rect 16865 5593 16899 5627
rect 17233 5593 17267 5627
rect 18061 5593 18095 5627
rect 22201 5593 22235 5627
rect 23949 5593 23983 5627
rect 1501 5525 1535 5559
rect 6745 5525 6779 5559
rect 9597 5525 9631 5559
rect 10701 5525 10735 5559
rect 12541 5525 12575 5559
rect 13737 5525 13771 5559
rect 17601 5525 17635 5559
rect 18521 5525 18555 5559
rect 19625 5525 19659 5559
rect 24409 5525 24443 5559
rect 24869 5525 24903 5559
rect 9321 5321 9355 5355
rect 9689 5321 9723 5355
rect 11529 5321 11563 5355
rect 12357 5321 12391 5355
rect 18061 5321 18095 5355
rect 19625 5321 19659 5355
rect 22753 5321 22787 5355
rect 9873 5253 9907 5287
rect 10425 5253 10459 5287
rect 10793 5253 10827 5287
rect 13921 5253 13955 5287
rect 14381 5253 14415 5287
rect 19717 5253 19751 5287
rect 22293 5253 22327 5287
rect 22661 5253 22695 5287
rect 24032 5253 24066 5287
rect 7941 5185 7975 5219
rect 8208 5185 8242 5219
rect 9597 5185 9631 5219
rect 10149 5185 10183 5219
rect 10241 5185 10275 5219
rect 10701 5185 10735 5219
rect 10977 5185 11011 5219
rect 11805 5185 11839 5219
rect 12081 5185 12115 5219
rect 12725 5185 12759 5219
rect 13001 5185 13035 5219
rect 13645 5185 13679 5219
rect 14197 5185 14231 5219
rect 14473 5185 14507 5219
rect 15117 5185 15151 5219
rect 15669 5185 15703 5219
rect 16129 5185 16163 5219
rect 16681 5185 16715 5219
rect 16948 5185 16982 5219
rect 18337 5185 18371 5219
rect 18613 5185 18647 5219
rect 21925 5185 21959 5219
rect 22109 5185 22143 5219
rect 23121 5185 23155 5219
rect 23305 5185 23339 5219
rect 10425 5117 10459 5151
rect 12633 5117 12667 5151
rect 13093 5117 13127 5151
rect 13921 5117 13955 5151
rect 15025 5117 15059 5151
rect 16037 5117 16071 5151
rect 23765 5117 23799 5151
rect 9873 5049 9907 5083
rect 10977 5049 11011 5083
rect 11713 4981 11747 5015
rect 12541 4981 12575 5015
rect 13185 4981 13219 5015
rect 13369 4981 13403 5015
rect 13737 4981 13771 5015
rect 14197 4981 14231 5015
rect 14749 4981 14783 5015
rect 15761 4981 15795 5015
rect 16313 4981 16347 5015
rect 23121 4981 23155 5015
rect 25145 4981 25179 5015
rect 9873 4777 9907 4811
rect 13185 4777 13219 4811
rect 16497 4777 16531 4811
rect 18153 4777 18187 4811
rect 20361 4777 20395 4811
rect 21005 4777 21039 4811
rect 15209 4709 15243 4743
rect 22661 4709 22695 4743
rect 13277 4641 13311 4675
rect 14381 4641 14415 4675
rect 21833 4641 21867 4675
rect 9689 4573 9723 4607
rect 10425 4573 10459 4607
rect 10609 4573 10643 4607
rect 11069 4573 11103 4607
rect 11437 4573 11471 4607
rect 12449 4573 12483 4607
rect 12725 4573 12759 4607
rect 13185 4573 13219 4607
rect 14105 4573 14139 4607
rect 15577 4573 15611 4607
rect 16129 4573 16163 4607
rect 16497 4573 16531 4607
rect 18429 4573 18463 4607
rect 18705 4573 18739 4607
rect 19349 4573 19383 4607
rect 19441 4573 19475 4607
rect 19717 4573 19751 4607
rect 19809 4573 19843 4607
rect 20821 4573 20855 4607
rect 21097 4573 21131 4607
rect 21373 4573 21407 4607
rect 21557 4573 21591 4607
rect 21741 4573 21775 4607
rect 22661 4573 22695 4607
rect 22753 4573 22787 4607
rect 23305 4573 23339 4607
rect 28365 4573 28399 4607
rect 9505 4505 9539 4539
rect 11621 4505 11655 4539
rect 13461 4505 13495 4539
rect 15393 4505 15427 4539
rect 17785 4505 17819 4539
rect 17969 4505 18003 4539
rect 18797 4505 18831 4539
rect 19533 4505 19567 4539
rect 23029 4505 23063 4539
rect 13001 4437 13035 4471
rect 16681 4437 16715 4471
rect 19809 4437 19843 4471
rect 20637 4437 20671 4471
rect 22937 4437 22971 4471
rect 23397 4437 23431 4471
rect 9781 4233 9815 4267
rect 14013 4233 14047 4267
rect 19441 4233 19475 4267
rect 21465 4233 21499 4267
rect 13645 4165 13679 4199
rect 15126 4165 15160 4199
rect 16957 4165 16991 4199
rect 18981 4165 19015 4199
rect 20352 4165 20386 4199
rect 8401 4097 8435 4131
rect 8668 4097 8702 4131
rect 10241 4097 10275 4131
rect 10425 4097 10459 4131
rect 11805 4097 11839 4131
rect 12265 4097 12299 4131
rect 12403 4097 12437 4131
rect 12541 4097 12575 4131
rect 12633 4097 12667 4131
rect 13369 4097 13403 4131
rect 16681 4097 16715 4131
rect 16773 4097 16807 4131
rect 17233 4097 17267 4131
rect 17417 4097 17451 4131
rect 17693 4097 17727 4131
rect 17969 4097 18003 4131
rect 19257 4097 19291 4131
rect 20085 4097 20119 4131
rect 22017 4097 22051 4131
rect 23958 4097 23992 4131
rect 11713 4029 11747 4063
rect 13461 4029 13495 4063
rect 15393 4029 15427 4063
rect 17325 4029 17359 4063
rect 19073 4029 19107 4063
rect 21925 4029 21959 4063
rect 22385 4029 22419 4063
rect 24225 4029 24259 4063
rect 13185 3961 13219 3995
rect 22845 3961 22879 3995
rect 10241 3893 10275 3927
rect 10609 3893 10643 3927
rect 12081 3893 12115 3927
rect 13369 3893 13403 3927
rect 16957 3893 16991 3927
rect 18981 3893 19015 3927
rect 11805 3689 11839 3723
rect 17601 3689 17635 3723
rect 17877 3689 17911 3723
rect 18337 3689 18371 3723
rect 19533 3689 19567 3723
rect 19993 3689 20027 3723
rect 20361 3689 20395 3723
rect 12173 3621 12207 3655
rect 13737 3621 13771 3655
rect 12357 3553 12391 3587
rect 13185 3553 13219 3587
rect 18061 3553 18095 3587
rect 19395 3553 19429 3587
rect 20729 3553 20763 3587
rect 10885 3485 10919 3519
rect 11161 3485 11195 3519
rect 12081 3485 12115 3519
rect 12909 3485 12943 3519
rect 13001 3485 13035 3519
rect 13461 3485 13495 3519
rect 16221 3485 16255 3519
rect 17877 3485 17911 3519
rect 18153 3485 18187 3519
rect 19257 3485 19291 3519
rect 19717 3485 19751 3519
rect 19993 3485 20027 3519
rect 20085 3485 20119 3519
rect 20996 3485 21030 3519
rect 24409 3485 24443 3519
rect 11437 3417 11471 3451
rect 11621 3417 11655 3451
rect 12357 3417 12391 3451
rect 13737 3417 13771 3451
rect 16488 3417 16522 3451
rect 24654 3417 24688 3451
rect 10983 3349 11017 3383
rect 11069 3349 11103 3383
rect 13185 3349 13219 3383
rect 13553 3349 13587 3383
rect 19717 3349 19751 3383
rect 22109 3349 22143 3383
rect 25789 3349 25823 3383
rect 8217 3145 8251 3179
rect 13369 3145 13403 3179
rect 20361 3145 20395 3179
rect 7604 3077 7638 3111
rect 7849 3009 7883 3043
rect 11713 3009 11747 3043
rect 11969 3009 12003 3043
rect 14482 3009 14516 3043
rect 14749 3009 14783 3043
rect 18981 3009 19015 3043
rect 19248 3009 19282 3043
rect 28089 3009 28123 3043
rect 13093 2873 13127 2907
rect 1501 2805 1535 2839
rect 6469 2805 6503 2839
rect 28273 2805 28307 2839
rect 17049 2601 17083 2635
rect 20729 2601 20763 2635
rect 1869 2533 1903 2567
rect 27813 2533 27847 2567
rect 19533 2465 19567 2499
rect 2421 2397 2455 2431
rect 3801 2397 3835 2431
rect 6561 2397 6595 2431
rect 12357 2397 12391 2431
rect 19257 2397 19291 2431
rect 20913 2397 20947 2431
rect 21189 2397 21223 2431
rect 22293 2397 22327 2431
rect 25237 2397 25271 2431
rect 26985 2397 27019 2431
rect 1685 2329 1719 2363
rect 5365 2329 5399 2363
rect 5733 2329 5767 2363
rect 16313 2329 16347 2363
rect 16957 2329 16991 2363
rect 27997 2329 28031 2363
rect 2237 2261 2271 2295
rect 4997 2261 5031 2295
rect 18797 2261 18831 2295
rect 22109 2261 22143 2295
rect 25421 2261 25455 2295
rect 27537 2261 27571 2295
<< metal1 >>
rect 1104 27770 28888 27792
rect 1104 27718 5582 27770
rect 5634 27718 5646 27770
rect 5698 27718 5710 27770
rect 5762 27718 5774 27770
rect 5826 27718 5838 27770
rect 5890 27718 14846 27770
rect 14898 27718 14910 27770
rect 14962 27718 14974 27770
rect 15026 27718 15038 27770
rect 15090 27718 15102 27770
rect 15154 27718 24110 27770
rect 24162 27718 24174 27770
rect 24226 27718 24238 27770
rect 24290 27718 24302 27770
rect 24354 27718 24366 27770
rect 24418 27718 28888 27770
rect 1104 27696 28888 27718
rect 2406 27588 2412 27600
rect 2367 27560 2412 27588
rect 2406 27548 2412 27560
rect 2464 27548 2470 27600
rect 3970 27588 3976 27600
rect 3931 27560 3976 27588
rect 3970 27548 3976 27560
rect 4028 27548 4034 27600
rect 16482 27548 16488 27600
rect 16540 27588 16546 27600
rect 16761 27591 16819 27597
rect 16761 27588 16773 27591
rect 16540 27560 16773 27588
rect 16540 27548 16546 27560
rect 16761 27557 16773 27560
rect 16807 27557 16819 27591
rect 19426 27588 19432 27600
rect 19387 27560 19432 27588
rect 16761 27551 16819 27557
rect 19426 27548 19432 27560
rect 19484 27548 19490 27600
rect 21266 27548 21272 27600
rect 21324 27588 21330 27600
rect 21821 27591 21879 27597
rect 21821 27588 21833 27591
rect 21324 27560 21833 27588
rect 21324 27548 21330 27560
rect 21821 27557 21833 27560
rect 21867 27557 21879 27591
rect 22370 27588 22376 27600
rect 22331 27560 22376 27588
rect 21821 27551 21879 27557
rect 22370 27548 22376 27560
rect 22428 27548 22434 27600
rect 23934 27588 23940 27600
rect 23895 27560 23940 27588
rect 23934 27548 23940 27560
rect 23992 27548 23998 27600
rect 25498 27588 25504 27600
rect 25459 27560 25504 27588
rect 25498 27548 25504 27560
rect 25556 27548 25562 27600
rect 25866 27588 25872 27600
rect 25827 27560 25872 27588
rect 25866 27548 25872 27560
rect 25924 27548 25930 27600
rect 27801 27591 27859 27597
rect 27801 27557 27813 27591
rect 27847 27588 27859 27591
rect 27982 27588 27988 27600
rect 27847 27560 27988 27588
rect 27847 27557 27859 27560
rect 27801 27551 27859 27557
rect 27982 27548 27988 27560
rect 28040 27548 28046 27600
rect 28258 27588 28264 27600
rect 28219 27560 28264 27588
rect 28258 27548 28264 27560
rect 28316 27548 28322 27600
rect 1670 27452 1676 27464
rect 1631 27424 1676 27452
rect 1670 27412 1676 27424
rect 1728 27412 1734 27464
rect 2424 27452 2452 27548
rect 2777 27455 2835 27461
rect 2777 27452 2789 27455
rect 2424 27424 2789 27452
rect 2777 27421 2789 27424
rect 2823 27421 2835 27455
rect 10502 27452 10508 27464
rect 10463 27424 10508 27452
rect 2777 27415 2835 27421
rect 10502 27412 10508 27424
rect 10560 27452 10566 27464
rect 10965 27455 11023 27461
rect 10965 27452 10977 27455
rect 10560 27424 10977 27452
rect 10560 27412 10566 27424
rect 10965 27421 10977 27424
rect 11011 27421 11023 27455
rect 10965 27415 11023 27421
rect 16945 27455 17003 27461
rect 16945 27421 16957 27455
rect 16991 27452 17003 27455
rect 18322 27452 18328 27464
rect 16991 27424 18328 27452
rect 16991 27421 17003 27424
rect 16945 27415 17003 27421
rect 18322 27412 18328 27424
rect 18380 27412 18386 27464
rect 22388 27452 22416 27548
rect 22741 27455 22799 27461
rect 22741 27452 22753 27455
rect 22388 27424 22753 27452
rect 22741 27421 22753 27424
rect 22787 27421 22799 27455
rect 23952 27452 23980 27548
rect 24673 27455 24731 27461
rect 24673 27452 24685 27455
rect 23952 27424 24685 27452
rect 22741 27415 22799 27421
rect 24673 27421 24685 27424
rect 24719 27421 24731 27455
rect 24673 27415 24731 27421
rect 25130 27412 25136 27464
rect 25188 27452 25194 27464
rect 25317 27455 25375 27461
rect 25317 27452 25329 27455
rect 25188 27424 25329 27452
rect 25188 27412 25194 27424
rect 25317 27421 25329 27424
rect 25363 27421 25375 27455
rect 25317 27415 25375 27421
rect 28077 27455 28135 27461
rect 28077 27421 28089 27455
rect 28123 27421 28135 27455
rect 28077 27415 28135 27421
rect 3142 27384 3148 27396
rect 3103 27356 3148 27384
rect 3142 27344 3148 27356
rect 3200 27344 3206 27396
rect 10689 27387 10747 27393
rect 10689 27353 10701 27387
rect 10735 27384 10747 27387
rect 10778 27384 10784 27396
rect 10735 27356 10784 27384
rect 10735 27353 10747 27356
rect 10689 27347 10747 27353
rect 10778 27344 10784 27356
rect 10836 27344 10842 27396
rect 25038 27384 25044 27396
rect 24999 27356 25044 27384
rect 25038 27344 25044 27356
rect 25096 27344 25102 27396
rect 1762 27316 1768 27328
rect 1723 27288 1768 27316
rect 1762 27276 1768 27288
rect 1820 27276 1826 27328
rect 22830 27316 22836 27328
rect 22791 27288 22836 27316
rect 22830 27276 22836 27288
rect 22888 27276 22894 27328
rect 23474 27276 23480 27328
rect 23532 27316 23538 27328
rect 28092 27316 28120 27415
rect 23532 27288 28120 27316
rect 23532 27276 23538 27288
rect 1104 27226 28888 27248
rect 1104 27174 10214 27226
rect 10266 27174 10278 27226
rect 10330 27174 10342 27226
rect 10394 27174 10406 27226
rect 10458 27174 10470 27226
rect 10522 27174 19478 27226
rect 19530 27174 19542 27226
rect 19594 27174 19606 27226
rect 19658 27174 19670 27226
rect 19722 27174 19734 27226
rect 19786 27174 28888 27226
rect 1104 27152 28888 27174
rect 1670 27072 1676 27124
rect 1728 27112 1734 27124
rect 2317 27115 2375 27121
rect 2317 27112 2329 27115
rect 1728 27084 2329 27112
rect 1728 27072 1734 27084
rect 2317 27081 2329 27084
rect 2363 27081 2375 27115
rect 23474 27112 23480 27124
rect 23435 27084 23480 27112
rect 2317 27075 2375 27081
rect 23474 27072 23480 27084
rect 23532 27072 23538 27124
rect 25130 27112 25136 27124
rect 25091 27084 25136 27112
rect 25130 27072 25136 27084
rect 25188 27072 25194 27124
rect 27522 27072 27528 27124
rect 27580 27112 27586 27124
rect 28261 27115 28319 27121
rect 28261 27112 28273 27115
rect 27580 27084 28273 27112
rect 27580 27072 27586 27084
rect 28261 27081 28273 27084
rect 28307 27081 28319 27115
rect 28261 27075 28319 27081
rect 22112 27016 23796 27044
rect 1394 26976 1400 26988
rect 1355 26948 1400 26976
rect 1394 26936 1400 26948
rect 1452 26976 1458 26988
rect 1949 26979 2007 26985
rect 1949 26976 1961 26979
rect 1452 26948 1961 26976
rect 1452 26936 1458 26948
rect 1949 26945 1961 26948
rect 1995 26945 2007 26979
rect 1949 26939 2007 26945
rect 20898 26868 20904 26920
rect 20956 26908 20962 26920
rect 22112 26917 22140 27016
rect 22370 26985 22376 26988
rect 22364 26939 22376 26985
rect 22428 26976 22434 26988
rect 23768 26985 23796 27016
rect 24026 26985 24032 26988
rect 23753 26979 23811 26985
rect 22428 26948 22464 26976
rect 22370 26936 22376 26939
rect 22428 26936 22434 26948
rect 23753 26945 23765 26979
rect 23799 26945 23811 26979
rect 23753 26939 23811 26945
rect 24020 26939 24032 26985
rect 24084 26976 24090 26988
rect 28074 26976 28080 26988
rect 24084 26948 24120 26976
rect 28035 26948 28080 26976
rect 24026 26936 24032 26939
rect 24084 26936 24090 26948
rect 28074 26936 28080 26948
rect 28132 26936 28138 26988
rect 22097 26911 22155 26917
rect 22097 26908 22109 26911
rect 20956 26880 22109 26908
rect 20956 26868 20962 26880
rect 22097 26877 22109 26880
rect 22143 26877 22155 26911
rect 22097 26871 22155 26877
rect 1578 26772 1584 26784
rect 1539 26744 1584 26772
rect 1578 26732 1584 26744
rect 1636 26732 1642 26784
rect 1104 26682 28888 26704
rect 1104 26630 5582 26682
rect 5634 26630 5646 26682
rect 5698 26630 5710 26682
rect 5762 26630 5774 26682
rect 5826 26630 5838 26682
rect 5890 26630 14846 26682
rect 14898 26630 14910 26682
rect 14962 26630 14974 26682
rect 15026 26630 15038 26682
rect 15090 26630 15102 26682
rect 15154 26630 24110 26682
rect 24162 26630 24174 26682
rect 24226 26630 24238 26682
rect 24290 26630 24302 26682
rect 24354 26630 24366 26682
rect 24418 26630 28888 26682
rect 1104 26608 28888 26630
rect 28350 26568 28356 26580
rect 28311 26540 28356 26568
rect 28350 26528 28356 26540
rect 28408 26528 28414 26580
rect 1394 26364 1400 26376
rect 1355 26336 1400 26364
rect 1394 26324 1400 26336
rect 1452 26324 1458 26376
rect 1104 26138 28888 26160
rect 1104 26086 10214 26138
rect 10266 26086 10278 26138
rect 10330 26086 10342 26138
rect 10394 26086 10406 26138
rect 10458 26086 10470 26138
rect 10522 26086 19478 26138
rect 19530 26086 19542 26138
rect 19594 26086 19606 26138
rect 19658 26086 19670 26138
rect 19722 26086 19734 26138
rect 19786 26086 28888 26138
rect 1104 26064 28888 26086
rect 1104 25594 28888 25616
rect 1104 25542 5582 25594
rect 5634 25542 5646 25594
rect 5698 25542 5710 25594
rect 5762 25542 5774 25594
rect 5826 25542 5838 25594
rect 5890 25542 14846 25594
rect 14898 25542 14910 25594
rect 14962 25542 14974 25594
rect 15026 25542 15038 25594
rect 15090 25542 15102 25594
rect 15154 25542 24110 25594
rect 24162 25542 24174 25594
rect 24226 25542 24238 25594
rect 24290 25542 24302 25594
rect 24354 25542 24366 25594
rect 24418 25542 28888 25594
rect 1104 25520 28888 25542
rect 27801 25279 27859 25285
rect 27801 25245 27813 25279
rect 27847 25276 27859 25279
rect 28350 25276 28356 25288
rect 27847 25248 28356 25276
rect 27847 25245 27859 25248
rect 27801 25239 27859 25245
rect 28350 25236 28356 25248
rect 28408 25236 28414 25288
rect 28166 25140 28172 25152
rect 28127 25112 28172 25140
rect 28166 25100 28172 25112
rect 28224 25100 28230 25152
rect 1104 25050 28888 25072
rect 1104 24998 10214 25050
rect 10266 24998 10278 25050
rect 10330 24998 10342 25050
rect 10394 24998 10406 25050
rect 10458 24998 10470 25050
rect 10522 24998 19478 25050
rect 19530 24998 19542 25050
rect 19594 24998 19606 25050
rect 19658 24998 19670 25050
rect 19722 24998 19734 25050
rect 19786 24998 28888 25050
rect 1104 24976 28888 24998
rect 9030 24828 9036 24880
rect 9088 24868 9094 24880
rect 12158 24868 12164 24880
rect 9088 24840 12164 24868
rect 9088 24828 9094 24840
rect 12158 24828 12164 24840
rect 12216 24828 12222 24880
rect 1394 24800 1400 24812
rect 1355 24772 1400 24800
rect 1394 24760 1400 24772
rect 1452 24800 1458 24812
rect 1949 24803 2007 24809
rect 1949 24800 1961 24803
rect 1452 24772 1961 24800
rect 1452 24760 1458 24772
rect 1949 24769 1961 24772
rect 1995 24769 2007 24803
rect 1949 24763 2007 24769
rect 14734 24760 14740 24812
rect 14792 24800 14798 24812
rect 14921 24803 14979 24809
rect 14921 24800 14933 24803
rect 14792 24772 14933 24800
rect 14792 24760 14798 24772
rect 14921 24769 14933 24772
rect 14967 24769 14979 24803
rect 14921 24763 14979 24769
rect 1581 24599 1639 24605
rect 1581 24565 1593 24599
rect 1627 24596 1639 24599
rect 1670 24596 1676 24608
rect 1627 24568 1676 24596
rect 1627 24565 1639 24568
rect 1581 24559 1639 24565
rect 1670 24556 1676 24568
rect 1728 24556 1734 24608
rect 14642 24556 14648 24608
rect 14700 24596 14706 24608
rect 14737 24599 14795 24605
rect 14737 24596 14749 24599
rect 14700 24568 14749 24596
rect 14700 24556 14706 24568
rect 14737 24565 14749 24568
rect 14783 24565 14795 24599
rect 14737 24559 14795 24565
rect 1104 24506 28888 24528
rect 1104 24454 5582 24506
rect 5634 24454 5646 24506
rect 5698 24454 5710 24506
rect 5762 24454 5774 24506
rect 5826 24454 5838 24506
rect 5890 24454 14846 24506
rect 14898 24454 14910 24506
rect 14962 24454 14974 24506
rect 15026 24454 15038 24506
rect 15090 24454 15102 24506
rect 15154 24454 24110 24506
rect 24162 24454 24174 24506
rect 24226 24454 24238 24506
rect 24290 24454 24302 24506
rect 24354 24454 24366 24506
rect 24418 24454 28888 24506
rect 1104 24432 28888 24454
rect 12894 24148 12900 24200
rect 12952 24188 12958 24200
rect 14642 24197 14648 24200
rect 14369 24191 14427 24197
rect 14369 24188 14381 24191
rect 12952 24160 14381 24188
rect 12952 24148 12958 24160
rect 14369 24157 14381 24160
rect 14415 24157 14427 24191
rect 14636 24188 14648 24197
rect 14603 24160 14648 24188
rect 14369 24151 14427 24157
rect 14636 24151 14648 24160
rect 14642 24148 14648 24151
rect 14700 24148 14706 24200
rect 16298 24148 16304 24200
rect 16356 24188 16362 24200
rect 16669 24191 16727 24197
rect 16669 24188 16681 24191
rect 16356 24160 16681 24188
rect 16356 24148 16362 24160
rect 16669 24157 16681 24160
rect 16715 24157 16727 24191
rect 16669 24151 16727 24157
rect 15562 24012 15568 24064
rect 15620 24052 15626 24064
rect 15749 24055 15807 24061
rect 15749 24052 15761 24055
rect 15620 24024 15761 24052
rect 15620 24012 15626 24024
rect 15749 24021 15761 24024
rect 15795 24021 15807 24055
rect 15749 24015 15807 24021
rect 16117 24055 16175 24061
rect 16117 24021 16129 24055
rect 16163 24052 16175 24055
rect 16390 24052 16396 24064
rect 16163 24024 16396 24052
rect 16163 24021 16175 24024
rect 16117 24015 16175 24021
rect 16390 24012 16396 24024
rect 16448 24012 16454 24064
rect 16853 24055 16911 24061
rect 16853 24021 16865 24055
rect 16899 24052 16911 24055
rect 16942 24052 16948 24064
rect 16899 24024 16948 24052
rect 16899 24021 16911 24024
rect 16853 24015 16911 24021
rect 16942 24012 16948 24024
rect 17000 24012 17006 24064
rect 17218 24052 17224 24064
rect 17179 24024 17224 24052
rect 17218 24012 17224 24024
rect 17276 24012 17282 24064
rect 1104 23962 28888 23984
rect 1104 23910 10214 23962
rect 10266 23910 10278 23962
rect 10330 23910 10342 23962
rect 10394 23910 10406 23962
rect 10458 23910 10470 23962
rect 10522 23910 19478 23962
rect 19530 23910 19542 23962
rect 19594 23910 19606 23962
rect 19658 23910 19670 23962
rect 19722 23910 19734 23962
rect 19786 23910 28888 23962
rect 1104 23888 28888 23910
rect 14645 23851 14703 23857
rect 14645 23817 14657 23851
rect 14691 23848 14703 23851
rect 14734 23848 14740 23860
rect 14691 23820 14740 23848
rect 14691 23817 14703 23820
rect 14645 23811 14703 23817
rect 14734 23808 14740 23820
rect 14792 23808 14798 23860
rect 16298 23848 16304 23860
rect 16259 23820 16304 23848
rect 16298 23808 16304 23820
rect 16356 23808 16362 23860
rect 16390 23808 16396 23860
rect 16448 23848 16454 23860
rect 22830 23848 22836 23860
rect 16448 23820 22836 23848
rect 16448 23808 16454 23820
rect 22830 23808 22836 23820
rect 22888 23808 22894 23860
rect 15286 23780 15292 23792
rect 15199 23752 15292 23780
rect 15286 23740 15292 23752
rect 15344 23780 15350 23792
rect 16408 23780 16436 23808
rect 17126 23780 17132 23792
rect 15344 23752 16436 23780
rect 16684 23752 17132 23780
rect 15344 23740 15350 23752
rect 14461 23715 14519 23721
rect 14461 23681 14473 23715
rect 14507 23712 14519 23715
rect 15381 23715 15439 23721
rect 14507 23684 14964 23712
rect 14507 23681 14519 23684
rect 14461 23675 14519 23681
rect 14277 23647 14335 23653
rect 14277 23613 14289 23647
rect 14323 23613 14335 23647
rect 14277 23607 14335 23613
rect 1394 23508 1400 23520
rect 1355 23480 1400 23508
rect 1394 23468 1400 23480
rect 1452 23468 1458 23520
rect 14292 23508 14320 23607
rect 14936 23585 14964 23684
rect 15381 23681 15393 23715
rect 15427 23712 15439 23715
rect 15562 23712 15568 23724
rect 15427 23684 15568 23712
rect 15427 23681 15439 23684
rect 15381 23675 15439 23681
rect 15562 23672 15568 23684
rect 15620 23672 15626 23724
rect 16114 23712 16120 23724
rect 16075 23684 16120 23712
rect 16114 23672 16120 23684
rect 16172 23672 16178 23724
rect 15470 23644 15476 23656
rect 15431 23616 15476 23644
rect 15470 23604 15476 23616
rect 15528 23604 15534 23656
rect 16684 23653 16712 23752
rect 17126 23740 17132 23752
rect 17184 23740 17190 23792
rect 20898 23780 20904 23792
rect 19352 23752 20760 23780
rect 20859 23752 20904 23780
rect 16942 23721 16948 23724
rect 16936 23712 16948 23721
rect 16903 23684 16948 23712
rect 16936 23675 16948 23684
rect 16942 23672 16948 23675
rect 17000 23672 17006 23724
rect 15933 23647 15991 23653
rect 15933 23613 15945 23647
rect 15979 23613 15991 23647
rect 15933 23607 15991 23613
rect 16669 23647 16727 23653
rect 16669 23613 16681 23647
rect 16715 23613 16727 23647
rect 16669 23607 16727 23613
rect 14921 23579 14979 23585
rect 14921 23545 14933 23579
rect 14967 23545 14979 23579
rect 14921 23539 14979 23545
rect 15654 23508 15660 23520
rect 14292 23480 15660 23508
rect 15654 23468 15660 23480
rect 15712 23508 15718 23520
rect 15948 23508 15976 23607
rect 19242 23536 19248 23588
rect 19300 23576 19306 23588
rect 19352 23585 19380 23752
rect 20732 23721 20760 23752
rect 20898 23740 20904 23752
rect 20956 23740 20962 23792
rect 19521 23715 19579 23721
rect 19521 23681 19533 23715
rect 19567 23712 19579 23715
rect 20717 23715 20775 23721
rect 19567 23684 20024 23712
rect 19567 23681 19579 23684
rect 19521 23675 19579 23681
rect 19337 23579 19395 23585
rect 19337 23576 19349 23579
rect 19300 23548 19349 23576
rect 19300 23536 19306 23548
rect 19337 23545 19349 23548
rect 19383 23545 19395 23579
rect 19337 23539 19395 23545
rect 15712 23480 15976 23508
rect 15712 23468 15718 23480
rect 17034 23468 17040 23520
rect 17092 23508 17098 23520
rect 19996 23517 20024 23684
rect 20717 23681 20729 23715
rect 20763 23681 20775 23715
rect 20717 23675 20775 23681
rect 18049 23511 18107 23517
rect 18049 23508 18061 23511
rect 17092 23480 18061 23508
rect 17092 23468 17098 23480
rect 18049 23477 18061 23480
rect 18095 23477 18107 23511
rect 18049 23471 18107 23477
rect 19981 23511 20039 23517
rect 19981 23477 19993 23511
rect 20027 23508 20039 23511
rect 21174 23508 21180 23520
rect 20027 23480 21180 23508
rect 20027 23477 20039 23480
rect 19981 23471 20039 23477
rect 21174 23468 21180 23480
rect 21232 23468 21238 23520
rect 28350 23508 28356 23520
rect 28311 23480 28356 23508
rect 28350 23468 28356 23480
rect 28408 23468 28414 23520
rect 1104 23418 28888 23440
rect 1104 23366 5582 23418
rect 5634 23366 5646 23418
rect 5698 23366 5710 23418
rect 5762 23366 5774 23418
rect 5826 23366 5838 23418
rect 5890 23366 14846 23418
rect 14898 23366 14910 23418
rect 14962 23366 14974 23418
rect 15026 23366 15038 23418
rect 15090 23366 15102 23418
rect 15154 23366 24110 23418
rect 24162 23366 24174 23418
rect 24226 23366 24238 23418
rect 24290 23366 24302 23418
rect 24354 23366 24366 23418
rect 24418 23366 28888 23418
rect 1104 23344 28888 23366
rect 15286 23304 15292 23316
rect 15247 23276 15292 23304
rect 15286 23264 15292 23276
rect 15344 23264 15350 23316
rect 16114 23264 16120 23316
rect 16172 23304 16178 23316
rect 16209 23307 16267 23313
rect 16209 23304 16221 23307
rect 16172 23276 16221 23304
rect 16172 23264 16178 23276
rect 16209 23273 16221 23276
rect 16255 23273 16267 23307
rect 16209 23267 16267 23273
rect 17218 23264 17224 23316
rect 17276 23304 17282 23316
rect 20530 23304 20536 23316
rect 17276 23276 20536 23304
rect 17276 23264 17282 23276
rect 20530 23264 20536 23276
rect 20588 23264 20594 23316
rect 15470 23196 15476 23248
rect 15528 23236 15534 23248
rect 16482 23236 16488 23248
rect 15528 23208 16488 23236
rect 15528 23196 15534 23208
rect 16482 23196 16488 23208
rect 16540 23236 16546 23248
rect 16540 23208 16804 23236
rect 16540 23196 16546 23208
rect 15565 23171 15623 23177
rect 15565 23137 15577 23171
rect 15611 23168 15623 23171
rect 15654 23168 15660 23180
rect 15611 23140 15660 23168
rect 15611 23137 15623 23140
rect 15565 23131 15623 23137
rect 15654 23128 15660 23140
rect 15712 23128 15718 23180
rect 16776 23177 16804 23208
rect 16761 23171 16819 23177
rect 16761 23137 16773 23171
rect 16807 23137 16819 23171
rect 16761 23131 16819 23137
rect 12618 23060 12624 23112
rect 12676 23100 12682 23112
rect 12805 23103 12863 23109
rect 12805 23100 12817 23103
rect 12676 23072 12817 23100
rect 12676 23060 12682 23072
rect 12805 23069 12817 23072
rect 12851 23069 12863 23103
rect 13446 23100 13452 23112
rect 13407 23072 13452 23100
rect 12805 23063 12863 23069
rect 13446 23060 13452 23072
rect 13504 23060 13510 23112
rect 15746 23100 15752 23112
rect 15707 23072 15752 23100
rect 15746 23060 15752 23072
rect 15804 23060 15810 23112
rect 16577 23103 16635 23109
rect 16577 23069 16589 23103
rect 16623 23096 16635 23103
rect 17218 23100 17224 23112
rect 16684 23096 17224 23100
rect 16623 23072 17224 23096
rect 16623 23069 16712 23072
rect 16577 23068 16712 23069
rect 16577 23063 16635 23068
rect 17218 23060 17224 23072
rect 17276 23060 17282 23112
rect 17773 23103 17831 23109
rect 17773 23100 17785 23103
rect 17328 23072 17785 23100
rect 15933 23035 15991 23041
rect 15933 23001 15945 23035
rect 15979 23032 15991 23035
rect 17328 23032 17356 23072
rect 17773 23069 17785 23072
rect 17819 23069 17831 23103
rect 18414 23100 18420 23112
rect 18375 23072 18420 23100
rect 17773 23063 17831 23069
rect 18414 23060 18420 23072
rect 18472 23060 18478 23112
rect 18874 23100 18880 23112
rect 18835 23072 18880 23100
rect 18874 23060 18880 23072
rect 18932 23060 18938 23112
rect 19978 23060 19984 23112
rect 20036 23100 20042 23112
rect 20073 23103 20131 23109
rect 20073 23100 20085 23103
rect 20036 23072 20085 23100
rect 20036 23060 20042 23072
rect 20073 23069 20085 23072
rect 20119 23069 20131 23103
rect 20254 23100 20260 23112
rect 20215 23072 20260 23100
rect 20073 23063 20131 23069
rect 20254 23060 20260 23072
rect 20312 23060 20318 23112
rect 15979 23004 17356 23032
rect 17405 23035 17463 23041
rect 15979 23001 15991 23004
rect 15933 22995 15991 23001
rect 17405 23001 17417 23035
rect 17451 23032 17463 23035
rect 19242 23032 19248 23044
rect 17451 23004 19248 23032
rect 17451 23001 17463 23004
rect 17405 22995 17463 23001
rect 19242 22992 19248 23004
rect 19300 22992 19306 23044
rect 19334 22992 19340 23044
rect 19392 23032 19398 23044
rect 19521 23035 19579 23041
rect 19521 23032 19533 23035
rect 19392 23004 19533 23032
rect 19392 22992 19398 23004
rect 19521 23001 19533 23004
rect 19567 23001 19579 23035
rect 19521 22995 19579 23001
rect 19705 23035 19763 23041
rect 19705 23001 19717 23035
rect 19751 23032 19763 23035
rect 19886 23032 19892 23044
rect 19751 23004 19892 23032
rect 19751 23001 19763 23004
rect 19705 22995 19763 23001
rect 19886 22992 19892 23004
rect 19944 22992 19950 23044
rect 12986 22964 12992 22976
rect 12947 22936 12992 22964
rect 12986 22924 12992 22936
rect 13044 22924 13050 22976
rect 13262 22964 13268 22976
rect 13223 22936 13268 22964
rect 13262 22924 13268 22936
rect 13320 22924 13326 22976
rect 15562 22924 15568 22976
rect 15620 22964 15626 22976
rect 15838 22964 15844 22976
rect 15620 22936 15844 22964
rect 15620 22924 15626 22936
rect 15838 22924 15844 22936
rect 15896 22924 15902 22976
rect 16669 22967 16727 22973
rect 16669 22933 16681 22967
rect 16715 22964 16727 22967
rect 17034 22964 17040 22976
rect 16715 22936 17040 22964
rect 16715 22933 16727 22936
rect 16669 22927 16727 22933
rect 17034 22924 17040 22936
rect 17092 22924 17098 22976
rect 17126 22924 17132 22976
rect 17184 22964 17190 22976
rect 17313 22967 17371 22973
rect 17313 22964 17325 22967
rect 17184 22936 17325 22964
rect 17184 22924 17190 22936
rect 17313 22933 17325 22936
rect 17359 22933 17371 22967
rect 17954 22964 17960 22976
rect 17915 22936 17960 22964
rect 17313 22927 17371 22933
rect 17954 22924 17960 22936
rect 18012 22924 18018 22976
rect 18230 22964 18236 22976
rect 18191 22936 18236 22964
rect 18230 22924 18236 22936
rect 18288 22924 18294 22976
rect 18690 22964 18696 22976
rect 18651 22936 18696 22964
rect 18690 22924 18696 22936
rect 18748 22924 18754 22976
rect 20441 22967 20499 22973
rect 20441 22933 20453 22967
rect 20487 22964 20499 22967
rect 21450 22964 21456 22976
rect 20487 22936 21456 22964
rect 20487 22933 20499 22936
rect 20441 22927 20499 22933
rect 21450 22924 21456 22936
rect 21508 22924 21514 22976
rect 1104 22874 28888 22896
rect 1104 22822 10214 22874
rect 10266 22822 10278 22874
rect 10330 22822 10342 22874
rect 10394 22822 10406 22874
rect 10458 22822 10470 22874
rect 10522 22822 19478 22874
rect 19530 22822 19542 22874
rect 19594 22822 19606 22874
rect 19658 22822 19670 22874
rect 19722 22822 19734 22874
rect 19786 22822 28888 22874
rect 1104 22800 28888 22822
rect 12618 22760 12624 22772
rect 12579 22732 12624 22760
rect 12618 22720 12624 22732
rect 12676 22720 12682 22772
rect 14277 22763 14335 22769
rect 14277 22729 14289 22763
rect 14323 22760 14335 22763
rect 15013 22763 15071 22769
rect 15013 22760 15025 22763
rect 14323 22732 15025 22760
rect 14323 22729 14335 22732
rect 14277 22723 14335 22729
rect 15013 22729 15025 22732
rect 15059 22760 15071 22763
rect 15838 22760 15844 22772
rect 15059 22732 15608 22760
rect 15059 22729 15071 22732
rect 15013 22723 15071 22729
rect 12526 22692 12532 22704
rect 12360 22664 12532 22692
rect 10870 22584 10876 22636
rect 10928 22624 10934 22636
rect 12360 22633 12388 22664
rect 12526 22652 12532 22664
rect 12584 22652 12590 22704
rect 12986 22652 12992 22704
rect 13044 22692 13050 22704
rect 13142 22695 13200 22701
rect 13142 22692 13154 22695
rect 13044 22664 13154 22692
rect 13044 22652 13050 22664
rect 13142 22661 13154 22664
rect 13188 22661 13200 22695
rect 13142 22655 13200 22661
rect 14921 22695 14979 22701
rect 14921 22661 14933 22695
rect 14967 22692 14979 22695
rect 15286 22692 15292 22704
rect 14967 22664 15292 22692
rect 14967 22661 14979 22664
rect 14921 22655 14979 22661
rect 15286 22652 15292 22664
rect 15344 22652 15350 22704
rect 12345 22627 12403 22633
rect 12345 22624 12357 22627
rect 10928 22596 12357 22624
rect 10928 22584 10934 22596
rect 12345 22593 12357 22596
rect 12391 22593 12403 22627
rect 12345 22587 12403 22593
rect 12437 22627 12495 22633
rect 12437 22593 12449 22627
rect 12483 22593 12495 22627
rect 12894 22624 12900 22636
rect 12855 22596 12900 22624
rect 12437 22587 12495 22593
rect 10502 22420 10508 22432
rect 10463 22392 10508 22420
rect 10502 22380 10508 22392
rect 10560 22380 10566 22432
rect 12452 22420 12480 22587
rect 12894 22584 12900 22596
rect 12952 22584 12958 22636
rect 15580 22633 15608 22732
rect 15764 22732 15844 22760
rect 15764 22701 15792 22732
rect 15838 22720 15844 22732
rect 15896 22720 15902 22772
rect 16117 22763 16175 22769
rect 16117 22729 16129 22763
rect 16163 22760 16175 22763
rect 17218 22760 17224 22772
rect 16163 22732 17224 22760
rect 16163 22729 16175 22732
rect 16117 22723 16175 22729
rect 17218 22720 17224 22732
rect 17276 22720 17282 22772
rect 15749 22695 15807 22701
rect 15749 22661 15761 22695
rect 15795 22661 15807 22695
rect 15749 22655 15807 22661
rect 17126 22652 17132 22704
rect 17184 22692 17190 22704
rect 18592 22695 18650 22701
rect 17184 22664 18092 22692
rect 17184 22652 17190 22664
rect 15565 22627 15623 22633
rect 15565 22593 15577 22627
rect 15611 22593 15623 22627
rect 15838 22624 15844 22636
rect 15799 22596 15844 22624
rect 15565 22587 15623 22593
rect 15838 22584 15844 22596
rect 15896 22584 15902 22636
rect 15930 22584 15936 22636
rect 15988 22624 15994 22636
rect 17793 22627 17851 22633
rect 15988 22596 16033 22624
rect 15988 22584 15994 22596
rect 17793 22593 17805 22627
rect 17839 22624 17851 22627
rect 17954 22624 17960 22636
rect 17839 22596 17960 22624
rect 17839 22593 17851 22596
rect 17793 22587 17851 22593
rect 17954 22584 17960 22596
rect 18012 22584 18018 22636
rect 18064 22633 18092 22664
rect 18592 22661 18604 22695
rect 18638 22692 18650 22695
rect 18690 22692 18696 22704
rect 18638 22664 18696 22692
rect 18638 22661 18650 22664
rect 18592 22655 18650 22661
rect 18690 22652 18696 22664
rect 18748 22652 18754 22704
rect 20898 22652 20904 22704
rect 20956 22692 20962 22704
rect 20956 22664 21496 22692
rect 20956 22652 20962 22664
rect 18049 22627 18107 22633
rect 18049 22593 18061 22627
rect 18095 22624 18107 22627
rect 18325 22627 18383 22633
rect 18325 22624 18337 22627
rect 18095 22596 18337 22624
rect 18095 22593 18107 22596
rect 18049 22587 18107 22593
rect 18325 22593 18337 22596
rect 18371 22593 18383 22627
rect 19334 22624 19340 22636
rect 18325 22587 18383 22593
rect 18432 22596 19340 22624
rect 14182 22516 14188 22568
rect 14240 22556 14246 22568
rect 15105 22559 15163 22565
rect 15105 22556 15117 22559
rect 14240 22528 15117 22556
rect 14240 22516 14246 22528
rect 15105 22525 15117 22528
rect 15151 22556 15163 22559
rect 18432 22556 18460 22596
rect 19334 22584 19340 22596
rect 19392 22624 19398 22636
rect 20622 22624 20628 22636
rect 19392 22596 20628 22624
rect 19392 22584 19398 22596
rect 20622 22584 20628 22596
rect 20680 22584 20686 22636
rect 21197 22627 21255 22633
rect 21197 22593 21209 22627
rect 21243 22624 21255 22627
rect 21358 22624 21364 22636
rect 21243 22596 21364 22624
rect 21243 22593 21255 22596
rect 21197 22587 21255 22593
rect 21358 22584 21364 22596
rect 21416 22584 21422 22636
rect 21468 22633 21496 22664
rect 21453 22627 21511 22633
rect 21453 22593 21465 22627
rect 21499 22593 21511 22627
rect 21453 22587 21511 22593
rect 15151 22528 16574 22556
rect 15151 22525 15163 22528
rect 15105 22519 15163 22525
rect 13906 22448 13912 22500
rect 13964 22488 13970 22500
rect 15838 22488 15844 22500
rect 13964 22460 15844 22488
rect 13964 22448 13970 22460
rect 15838 22448 15844 22460
rect 15896 22448 15902 22500
rect 16546 22488 16574 22528
rect 18340 22528 18460 22556
rect 16546 22460 17172 22488
rect 14553 22423 14611 22429
rect 14553 22420 14565 22423
rect 12452 22392 14565 22420
rect 14553 22389 14565 22392
rect 14599 22389 14611 22423
rect 16666 22420 16672 22432
rect 16627 22392 16672 22420
rect 14553 22383 14611 22389
rect 16666 22380 16672 22392
rect 16724 22380 16730 22432
rect 17144 22420 17172 22460
rect 18340 22420 18368 22528
rect 20073 22491 20131 22497
rect 20073 22488 20085 22491
rect 19536 22460 20085 22488
rect 17144 22392 18368 22420
rect 19058 22380 19064 22432
rect 19116 22420 19122 22432
rect 19536 22420 19564 22460
rect 20073 22457 20085 22460
rect 20119 22457 20131 22491
rect 20073 22451 20131 22457
rect 19702 22420 19708 22432
rect 19116 22392 19564 22420
rect 19663 22392 19708 22420
rect 19116 22380 19122 22392
rect 19702 22380 19708 22392
rect 19760 22380 19766 22432
rect 1104 22330 28888 22352
rect 1104 22278 5582 22330
rect 5634 22278 5646 22330
rect 5698 22278 5710 22330
rect 5762 22278 5774 22330
rect 5826 22278 5838 22330
rect 5890 22278 14846 22330
rect 14898 22278 14910 22330
rect 14962 22278 14974 22330
rect 15026 22278 15038 22330
rect 15090 22278 15102 22330
rect 15154 22278 24110 22330
rect 24162 22278 24174 22330
rect 24226 22278 24238 22330
rect 24290 22278 24302 22330
rect 24354 22278 24366 22330
rect 24418 22278 28888 22330
rect 1104 22256 28888 22278
rect 15746 22176 15752 22228
rect 15804 22216 15810 22228
rect 16209 22219 16267 22225
rect 16209 22216 16221 22219
rect 15804 22188 16221 22216
rect 15804 22176 15810 22188
rect 16209 22185 16221 22188
rect 16255 22185 16267 22219
rect 16209 22179 16267 22185
rect 16666 22176 16672 22228
rect 16724 22216 16730 22228
rect 17586 22216 17592 22228
rect 16724 22188 17592 22216
rect 16724 22176 16730 22188
rect 17586 22176 17592 22188
rect 17644 22176 17650 22228
rect 18874 22216 18880 22228
rect 18835 22188 18880 22216
rect 18874 22176 18880 22188
rect 18932 22176 18938 22228
rect 20254 22216 20260 22228
rect 20215 22188 20260 22216
rect 20254 22176 20260 22188
rect 20312 22176 20318 22228
rect 21269 22219 21327 22225
rect 21269 22185 21281 22219
rect 21315 22216 21327 22219
rect 21358 22216 21364 22228
rect 21315 22188 21364 22216
rect 21315 22185 21327 22188
rect 21269 22179 21327 22185
rect 21358 22176 21364 22188
rect 21416 22176 21422 22228
rect 16482 22108 16488 22160
rect 16540 22148 16546 22160
rect 18782 22148 18788 22160
rect 16540 22120 16804 22148
rect 16540 22108 16546 22120
rect 16298 22040 16304 22092
rect 16356 22080 16362 22092
rect 16500 22080 16528 22108
rect 16776 22094 16804 22120
rect 17476 22120 18788 22148
rect 16776 22089 16841 22094
rect 16356 22052 16528 22080
rect 16761 22083 16841 22089
rect 16356 22040 16362 22052
rect 16761 22049 16773 22083
rect 16807 22066 16841 22083
rect 16807 22049 16819 22066
rect 16761 22043 16819 22049
rect 7558 21972 7564 22024
rect 7616 22012 7622 22024
rect 7837 22015 7895 22021
rect 7837 22012 7849 22015
rect 7616 21984 7849 22012
rect 7616 21972 7622 21984
rect 7837 21981 7849 21984
rect 7883 21981 7895 22015
rect 7837 21975 7895 21981
rect 9585 22015 9643 22021
rect 9585 21981 9597 22015
rect 9631 22012 9643 22015
rect 9674 22012 9680 22024
rect 9631 21984 9680 22012
rect 9631 21981 9643 21984
rect 9585 21975 9643 21981
rect 9674 21972 9680 21984
rect 9732 21972 9738 22024
rect 10321 22015 10379 22021
rect 10321 21981 10333 22015
rect 10367 22012 10379 22015
rect 10502 22012 10508 22024
rect 10367 21984 10508 22012
rect 10367 21981 10379 21984
rect 10321 21975 10379 21981
rect 10502 21972 10508 21984
rect 10560 21972 10566 22024
rect 12069 22015 12127 22021
rect 12069 21981 12081 22015
rect 12115 22012 12127 22015
rect 12345 22015 12403 22021
rect 12345 22012 12357 22015
rect 12115 21984 12357 22012
rect 12115 21981 12127 21984
rect 12069 21975 12127 21981
rect 12345 21981 12357 21984
rect 12391 22012 12403 22015
rect 12434 22012 12440 22024
rect 12391 21984 12440 22012
rect 12391 21981 12403 21984
rect 12345 21975 12403 21981
rect 12434 21972 12440 21984
rect 12492 22012 12498 22024
rect 12894 22012 12900 22024
rect 12492 21984 12900 22012
rect 12492 21972 12498 21984
rect 12894 21972 12900 21984
rect 12952 21972 12958 22024
rect 15657 22015 15715 22021
rect 15657 21981 15669 22015
rect 15703 22012 15715 22015
rect 17126 22012 17132 22024
rect 15703 21984 17132 22012
rect 15703 21981 15715 21984
rect 15657 21975 15715 21981
rect 17126 21972 17132 21984
rect 17184 21972 17190 22024
rect 17218 21972 17224 22024
rect 17276 22012 17282 22024
rect 17476 22021 17504 22120
rect 18782 22108 18788 22120
rect 18840 22108 18846 22160
rect 19058 22108 19064 22160
rect 19116 22148 19122 22160
rect 19116 22120 20760 22148
rect 19116 22108 19122 22120
rect 18966 22080 18972 22092
rect 17696 22052 18972 22080
rect 17586 22021 17592 22024
rect 17320 22015 17378 22021
rect 17320 22012 17332 22015
rect 17276 21984 17332 22012
rect 17276 21972 17282 21984
rect 17320 21981 17332 21984
rect 17366 21981 17378 22015
rect 17320 21975 17378 21981
rect 17451 22015 17509 22021
rect 17451 21981 17463 22015
rect 17497 21981 17509 22015
rect 17451 21975 17509 21981
rect 17543 22015 17592 22021
rect 17543 21981 17555 22015
rect 17589 21981 17592 22015
rect 17543 21975 17592 21981
rect 17586 21972 17592 21975
rect 17644 21972 17650 22024
rect 17696 22021 17724 22052
rect 18966 22040 18972 22052
rect 19024 22040 19030 22092
rect 19886 22080 19892 22092
rect 19847 22052 19892 22080
rect 19886 22040 19892 22052
rect 19944 22040 19950 22092
rect 20732 22089 20760 22120
rect 20717 22083 20775 22089
rect 20717 22049 20729 22083
rect 20763 22080 20775 22083
rect 20901 22083 20959 22089
rect 20763 22052 20797 22080
rect 20763 22049 20775 22052
rect 20717 22043 20775 22049
rect 20901 22049 20913 22083
rect 20947 22049 20959 22083
rect 20901 22043 20959 22049
rect 17678 22015 17736 22021
rect 17678 21981 17690 22015
rect 17724 21981 17736 22015
rect 17678 21975 17736 21981
rect 17778 22015 17836 22021
rect 17778 21981 17790 22015
rect 17824 21981 17836 22015
rect 18598 22012 18604 22024
rect 18559 21984 18604 22012
rect 17778 21975 17836 21981
rect 10134 21944 10140 21956
rect 10095 21916 10140 21944
rect 10134 21904 10140 21916
rect 10192 21904 10198 21956
rect 11606 21904 11612 21956
rect 11664 21944 11670 21956
rect 11802 21947 11860 21953
rect 11802 21944 11814 21947
rect 11664 21916 11814 21944
rect 11664 21904 11670 21916
rect 11802 21913 11814 21916
rect 11848 21913 11860 21947
rect 11802 21907 11860 21913
rect 12612 21947 12670 21953
rect 12612 21913 12624 21947
rect 12658 21944 12670 21947
rect 13262 21944 13268 21956
rect 12658 21916 13268 21944
rect 12658 21913 12670 21916
rect 12612 21907 12670 21913
rect 13262 21904 13268 21916
rect 13320 21904 13326 21956
rect 15412 21947 15470 21953
rect 15412 21913 15424 21947
rect 15458 21944 15470 21947
rect 16482 21944 16488 21956
rect 15458 21916 16488 21944
rect 15458 21913 15470 21916
rect 15412 21907 15470 21913
rect 16482 21904 16488 21916
rect 16540 21904 16546 21956
rect 7926 21836 7932 21888
rect 7984 21876 7990 21888
rect 8021 21879 8079 21885
rect 8021 21876 8033 21879
rect 7984 21848 8033 21876
rect 7984 21836 7990 21848
rect 8021 21845 8033 21848
rect 8067 21845 8079 21879
rect 9398 21876 9404 21888
rect 9359 21848 9404 21876
rect 8021 21839 8079 21845
rect 9398 21836 9404 21848
rect 9456 21836 9462 21888
rect 10689 21879 10747 21885
rect 10689 21845 10701 21879
rect 10735 21876 10747 21879
rect 12710 21876 12716 21888
rect 10735 21848 12716 21876
rect 10735 21845 10747 21848
rect 10689 21839 10747 21845
rect 12710 21836 12716 21848
rect 12768 21836 12774 21888
rect 13725 21879 13783 21885
rect 13725 21845 13737 21879
rect 13771 21876 13783 21879
rect 13906 21876 13912 21888
rect 13771 21848 13912 21876
rect 13771 21845 13783 21848
rect 13725 21839 13783 21845
rect 13906 21836 13912 21848
rect 13964 21836 13970 21888
rect 13998 21836 14004 21888
rect 14056 21876 14062 21888
rect 14277 21879 14335 21885
rect 14277 21876 14289 21879
rect 14056 21848 14289 21876
rect 14056 21836 14062 21848
rect 14277 21845 14289 21848
rect 14323 21845 14335 21879
rect 16574 21876 16580 21888
rect 16535 21848 16580 21876
rect 14277 21839 14335 21845
rect 16574 21836 16580 21848
rect 16632 21836 16638 21888
rect 16666 21836 16672 21888
rect 16724 21876 16730 21888
rect 16724 21848 16769 21876
rect 16724 21836 16730 21848
rect 17034 21836 17040 21888
rect 17092 21876 17098 21888
rect 17793 21876 17821 21975
rect 18598 21972 18604 21984
rect 18656 21972 18662 22024
rect 18690 21972 18696 22024
rect 18748 22012 18754 22024
rect 18748 21984 18793 22012
rect 18748 21972 18754 21984
rect 20530 21972 20536 22024
rect 20588 22012 20594 22024
rect 20625 22015 20683 22021
rect 20625 22012 20637 22015
rect 20588 21984 20637 22012
rect 20588 21972 20594 21984
rect 20625 21981 20637 21984
rect 20671 21981 20683 22015
rect 20625 21975 20683 21981
rect 18782 21904 18788 21956
rect 18840 21944 18846 21956
rect 19702 21944 19708 21956
rect 18840 21916 19708 21944
rect 18840 21904 18846 21916
rect 19702 21904 19708 21916
rect 19760 21904 19766 21956
rect 19886 21904 19892 21956
rect 19944 21944 19950 21956
rect 20916 21944 20944 22043
rect 21450 22012 21456 22024
rect 21411 21984 21456 22012
rect 21450 21972 21456 21984
rect 21508 21972 21514 22024
rect 19944 21916 20944 21944
rect 19944 21904 19950 21916
rect 17954 21876 17960 21888
rect 17092 21848 17821 21876
rect 17915 21848 17960 21876
rect 17092 21836 17098 21848
rect 17954 21836 17960 21848
rect 18012 21836 18018 21888
rect 18690 21836 18696 21888
rect 18748 21876 18754 21888
rect 19245 21879 19303 21885
rect 19245 21876 19257 21879
rect 18748 21848 19257 21876
rect 18748 21836 18754 21848
rect 19245 21845 19257 21848
rect 19291 21845 19303 21879
rect 19245 21839 19303 21845
rect 19334 21836 19340 21888
rect 19392 21876 19398 21888
rect 19613 21879 19671 21885
rect 19613 21876 19625 21879
rect 19392 21848 19625 21876
rect 19392 21836 19398 21848
rect 19613 21845 19625 21848
rect 19659 21876 19671 21879
rect 21729 21879 21787 21885
rect 21729 21876 21741 21879
rect 19659 21848 21741 21876
rect 19659 21845 19671 21848
rect 19613 21839 19671 21845
rect 21729 21845 21741 21848
rect 21775 21845 21787 21879
rect 21729 21839 21787 21845
rect 1104 21786 28888 21808
rect 1104 21734 10214 21786
rect 10266 21734 10278 21786
rect 10330 21734 10342 21786
rect 10394 21734 10406 21786
rect 10458 21734 10470 21786
rect 10522 21734 19478 21786
rect 19530 21734 19542 21786
rect 19594 21734 19606 21786
rect 19658 21734 19670 21786
rect 19722 21734 19734 21786
rect 19786 21734 28888 21786
rect 1104 21712 28888 21734
rect 9766 21632 9772 21684
rect 9824 21672 9830 21684
rect 10689 21675 10747 21681
rect 10689 21672 10701 21675
rect 9824 21644 10701 21672
rect 9824 21632 9830 21644
rect 10689 21641 10701 21644
rect 10735 21672 10747 21675
rect 11977 21675 12035 21681
rect 11977 21672 11989 21675
rect 10735 21644 11989 21672
rect 10735 21641 10747 21644
rect 10689 21635 10747 21641
rect 11977 21641 11989 21644
rect 12023 21641 12035 21675
rect 11977 21635 12035 21641
rect 12897 21675 12955 21681
rect 12897 21641 12909 21675
rect 12943 21672 12955 21675
rect 13446 21672 13452 21684
rect 12943 21644 13452 21672
rect 12943 21641 12955 21644
rect 12897 21635 12955 21641
rect 13446 21632 13452 21644
rect 13504 21632 13510 21684
rect 13906 21632 13912 21684
rect 13964 21672 13970 21684
rect 14001 21675 14059 21681
rect 14001 21672 14013 21675
rect 13964 21644 14013 21672
rect 13964 21632 13970 21644
rect 14001 21641 14013 21644
rect 14047 21641 14059 21675
rect 14001 21635 14059 21641
rect 16482 21632 16488 21684
rect 16540 21672 16546 21684
rect 16669 21675 16727 21681
rect 16669 21672 16681 21675
rect 16540 21644 16681 21672
rect 16540 21632 16546 21644
rect 16669 21641 16681 21644
rect 16715 21641 16727 21675
rect 16669 21635 16727 21641
rect 18414 21632 18420 21684
rect 18472 21672 18478 21684
rect 19153 21675 19211 21681
rect 19153 21672 19165 21675
rect 18472 21644 19165 21672
rect 18472 21632 18478 21644
rect 19153 21641 19165 21644
rect 19199 21641 19211 21675
rect 19153 21635 19211 21641
rect 20530 21632 20536 21684
rect 20588 21672 20594 21684
rect 21361 21675 21419 21681
rect 21361 21672 21373 21675
rect 20588 21644 21373 21672
rect 20588 21632 20594 21644
rect 21361 21641 21373 21644
rect 21407 21672 21419 21675
rect 25038 21672 25044 21684
rect 21407 21644 25044 21672
rect 21407 21641 21419 21644
rect 21361 21635 21419 21641
rect 25038 21632 25044 21644
rect 25096 21632 25102 21684
rect 7668 21576 9168 21604
rect 6822 21496 6828 21548
rect 6880 21536 6886 21548
rect 7668 21545 7696 21576
rect 7926 21545 7932 21548
rect 7653 21539 7711 21545
rect 7653 21536 7665 21539
rect 6880 21508 7665 21536
rect 6880 21496 6886 21508
rect 7653 21505 7665 21508
rect 7699 21505 7711 21539
rect 7920 21536 7932 21545
rect 7887 21508 7932 21536
rect 7653 21499 7711 21505
rect 7920 21499 7932 21508
rect 7926 21496 7932 21499
rect 7984 21496 7990 21548
rect 9140 21480 9168 21576
rect 9398 21564 9404 21616
rect 9456 21604 9462 21616
rect 9554 21607 9612 21613
rect 9554 21604 9566 21607
rect 9456 21576 9566 21604
rect 9456 21564 9462 21576
rect 9554 21573 9566 21576
rect 9600 21573 9612 21607
rect 9554 21567 9612 21573
rect 11885 21607 11943 21613
rect 11885 21573 11897 21607
rect 11931 21604 11943 21607
rect 12618 21604 12624 21616
rect 11931 21576 12624 21604
rect 11931 21573 11943 21576
rect 11885 21567 11943 21573
rect 12618 21564 12624 21576
rect 12676 21564 12682 21616
rect 15105 21607 15163 21613
rect 15105 21604 15117 21607
rect 13924 21576 15117 21604
rect 10965 21539 11023 21545
rect 10965 21505 10977 21539
rect 11011 21536 11023 21539
rect 11146 21536 11152 21548
rect 11011 21508 11152 21536
rect 11011 21505 11023 21508
rect 10965 21499 11023 21505
rect 11146 21496 11152 21508
rect 11204 21496 11210 21548
rect 13924 21545 13952 21576
rect 15105 21573 15117 21576
rect 15151 21573 15163 21607
rect 15105 21567 15163 21573
rect 15286 21564 15292 21616
rect 15344 21604 15350 21616
rect 17764 21607 17822 21613
rect 15344 21576 17724 21604
rect 15344 21564 15350 21576
rect 12713 21539 12771 21545
rect 12713 21505 12725 21539
rect 12759 21536 12771 21539
rect 13909 21539 13967 21545
rect 13909 21536 13921 21539
rect 12759 21508 13584 21536
rect 12759 21505 12771 21508
rect 12713 21499 12771 21505
rect 9122 21428 9128 21480
rect 9180 21468 9186 21480
rect 9309 21471 9367 21477
rect 9309 21468 9321 21471
rect 9180 21440 9321 21468
rect 9180 21428 9186 21440
rect 9309 21437 9321 21440
rect 9355 21437 9367 21471
rect 9309 21431 9367 21437
rect 12161 21471 12219 21477
rect 12161 21437 12173 21471
rect 12207 21468 12219 21471
rect 12342 21468 12348 21480
rect 12207 21440 12348 21468
rect 12207 21437 12219 21440
rect 12161 21431 12219 21437
rect 12342 21428 12348 21440
rect 12400 21428 12406 21480
rect 12526 21468 12532 21480
rect 12487 21440 12532 21468
rect 12526 21428 12532 21440
rect 12584 21428 12590 21480
rect 13556 21409 13584 21508
rect 13832 21508 13921 21536
rect 13541 21403 13599 21409
rect 8864 21372 9352 21400
rect 1394 21332 1400 21344
rect 1355 21304 1400 21332
rect 1394 21292 1400 21304
rect 1452 21292 1458 21344
rect 7650 21292 7656 21344
rect 7708 21332 7714 21344
rect 8864 21332 8892 21372
rect 9030 21332 9036 21344
rect 7708 21304 8892 21332
rect 8991 21304 9036 21332
rect 7708 21292 7714 21304
rect 9030 21292 9036 21304
rect 9088 21292 9094 21344
rect 9324 21332 9352 21372
rect 11072 21372 12434 21400
rect 11072 21332 11100 21372
rect 9324 21304 11100 21332
rect 11149 21335 11207 21341
rect 11149 21301 11161 21335
rect 11195 21332 11207 21335
rect 11330 21332 11336 21344
rect 11195 21304 11336 21332
rect 11195 21301 11207 21304
rect 11149 21295 11207 21301
rect 11330 21292 11336 21304
rect 11388 21292 11394 21344
rect 11514 21332 11520 21344
rect 11475 21304 11520 21332
rect 11514 21292 11520 21304
rect 11572 21292 11578 21344
rect 12406 21332 12434 21372
rect 13541 21369 13553 21403
rect 13587 21369 13599 21403
rect 13541 21363 13599 21369
rect 13265 21335 13323 21341
rect 13265 21332 13277 21335
rect 12406 21304 13277 21332
rect 13265 21301 13277 21304
rect 13311 21332 13323 21335
rect 13446 21332 13452 21344
rect 13311 21304 13452 21332
rect 13311 21301 13323 21304
rect 13265 21295 13323 21301
rect 13446 21292 13452 21304
rect 13504 21332 13510 21344
rect 13832 21332 13860 21508
rect 13909 21505 13921 21508
rect 13955 21505 13967 21539
rect 13909 21499 13967 21505
rect 13998 21496 14004 21548
rect 14056 21536 14062 21548
rect 15013 21539 15071 21545
rect 15013 21536 15025 21539
rect 14056 21508 15025 21536
rect 14056 21496 14062 21508
rect 15013 21505 15025 21508
rect 15059 21536 15071 21539
rect 15838 21536 15844 21548
rect 15059 21508 15844 21536
rect 15059 21505 15071 21508
rect 15013 21499 15071 21505
rect 15838 21496 15844 21508
rect 15896 21496 15902 21548
rect 15933 21539 15991 21545
rect 15933 21505 15945 21539
rect 15979 21505 15991 21539
rect 15933 21499 15991 21505
rect 16117 21539 16175 21545
rect 16117 21505 16129 21539
rect 16163 21536 16175 21539
rect 16853 21539 16911 21545
rect 16853 21536 16865 21539
rect 16163 21508 16865 21536
rect 16163 21505 16175 21508
rect 16117 21499 16175 21505
rect 16853 21505 16865 21508
rect 16899 21505 16911 21539
rect 16853 21499 16911 21505
rect 14182 21468 14188 21480
rect 14143 21440 14188 21468
rect 14182 21428 14188 21440
rect 14240 21428 14246 21480
rect 14921 21471 14979 21477
rect 14921 21437 14933 21471
rect 14967 21437 14979 21471
rect 15746 21468 15752 21480
rect 15707 21440 15752 21468
rect 14921 21431 14979 21437
rect 14936 21400 14964 21431
rect 15746 21428 15752 21440
rect 15804 21428 15810 21480
rect 15473 21403 15531 21409
rect 14936 21372 15056 21400
rect 13504 21304 13860 21332
rect 15028 21332 15056 21372
rect 15473 21369 15485 21403
rect 15519 21400 15531 21403
rect 15948 21400 15976 21499
rect 17126 21496 17132 21548
rect 17184 21536 17190 21548
rect 17497 21539 17555 21545
rect 17497 21536 17509 21539
rect 17184 21508 17509 21536
rect 17184 21496 17190 21508
rect 17497 21505 17509 21508
rect 17543 21505 17555 21539
rect 17696 21536 17724 21576
rect 17764 21573 17776 21607
rect 17810 21604 17822 21607
rect 18230 21604 18236 21616
rect 17810 21576 18236 21604
rect 17810 21573 17822 21576
rect 17764 21567 17822 21573
rect 18230 21564 18236 21576
rect 18288 21564 18294 21616
rect 18598 21564 18604 21616
rect 18656 21604 18662 21616
rect 18656 21576 19564 21604
rect 18656 21564 18662 21576
rect 17696 21508 18828 21536
rect 17497 21499 17555 21505
rect 15519 21372 15976 21400
rect 18800 21400 18828 21508
rect 18874 21496 18880 21548
rect 18932 21536 18938 21548
rect 19536 21545 19564 21576
rect 19337 21539 19395 21545
rect 19337 21536 19349 21539
rect 18932 21508 19349 21536
rect 18932 21496 18938 21508
rect 19337 21505 19349 21508
rect 19383 21505 19395 21539
rect 19337 21499 19395 21505
rect 19521 21539 19579 21545
rect 19521 21505 19533 21539
rect 19567 21536 19579 21539
rect 19610 21536 19616 21548
rect 19567 21508 19616 21536
rect 19567 21505 19579 21508
rect 19521 21499 19579 21505
rect 19610 21496 19616 21508
rect 19668 21536 19674 21548
rect 19978 21536 19984 21548
rect 19668 21508 19984 21536
rect 19668 21496 19674 21508
rect 19978 21496 19984 21508
rect 20036 21496 20042 21548
rect 20162 21536 20168 21548
rect 20123 21508 20168 21536
rect 20162 21496 20168 21508
rect 20220 21496 20226 21548
rect 20254 21496 20260 21548
rect 20312 21536 20318 21548
rect 20901 21539 20959 21545
rect 20901 21536 20913 21539
rect 20312 21508 20913 21536
rect 20312 21496 20318 21508
rect 20901 21505 20913 21508
rect 20947 21505 20959 21539
rect 20901 21499 20959 21505
rect 19978 21400 19984 21412
rect 18800 21372 19984 21400
rect 15519 21369 15531 21372
rect 15473 21363 15531 21369
rect 19978 21360 19984 21372
rect 20036 21360 20042 21412
rect 15562 21332 15568 21344
rect 15028 21304 15568 21332
rect 13504 21292 13510 21304
rect 15562 21292 15568 21304
rect 15620 21292 15626 21344
rect 16574 21292 16580 21344
rect 16632 21332 16638 21344
rect 17218 21332 17224 21344
rect 16632 21304 17224 21332
rect 16632 21292 16638 21304
rect 17218 21292 17224 21304
rect 17276 21292 17282 21344
rect 18414 21292 18420 21344
rect 18472 21332 18478 21344
rect 18877 21335 18935 21341
rect 18877 21332 18889 21335
rect 18472 21304 18889 21332
rect 18472 21292 18478 21304
rect 18877 21301 18889 21304
rect 18923 21301 18935 21335
rect 18877 21295 18935 21301
rect 20349 21335 20407 21341
rect 20349 21301 20361 21335
rect 20395 21332 20407 21335
rect 20898 21332 20904 21344
rect 20395 21304 20904 21332
rect 20395 21301 20407 21304
rect 20349 21295 20407 21301
rect 20898 21292 20904 21304
rect 20956 21292 20962 21344
rect 21085 21335 21143 21341
rect 21085 21301 21097 21335
rect 21131 21332 21143 21335
rect 21266 21332 21272 21344
rect 21131 21304 21272 21332
rect 21131 21301 21143 21304
rect 21085 21295 21143 21301
rect 21266 21292 21272 21304
rect 21324 21292 21330 21344
rect 1104 21242 28888 21264
rect 1104 21190 5582 21242
rect 5634 21190 5646 21242
rect 5698 21190 5710 21242
rect 5762 21190 5774 21242
rect 5826 21190 5838 21242
rect 5890 21190 14846 21242
rect 14898 21190 14910 21242
rect 14962 21190 14974 21242
rect 15026 21190 15038 21242
rect 15090 21190 15102 21242
rect 15154 21190 24110 21242
rect 24162 21190 24174 21242
rect 24226 21190 24238 21242
rect 24290 21190 24302 21242
rect 24354 21190 24366 21242
rect 24418 21190 28888 21242
rect 1104 21168 28888 21190
rect 7558 21128 7564 21140
rect 7519 21100 7564 21128
rect 7558 21088 7564 21100
rect 7616 21088 7622 21140
rect 11606 21128 11612 21140
rect 7760 21100 9444 21128
rect 11567 21100 11612 21128
rect 3142 21020 3148 21072
rect 3200 21060 3206 21072
rect 7650 21060 7656 21072
rect 3200 21032 7656 21060
rect 3200 21020 3206 21032
rect 7650 21020 7656 21032
rect 7708 21020 7714 21072
rect 6917 20995 6975 21001
rect 6917 20961 6929 20995
rect 6963 20992 6975 20995
rect 7193 20995 7251 21001
rect 7193 20992 7205 20995
rect 6963 20964 7205 20992
rect 6963 20961 6975 20964
rect 6917 20955 6975 20961
rect 7193 20961 7205 20964
rect 7239 20992 7251 20995
rect 7760 20992 7788 21100
rect 9416 21072 9444 21100
rect 11606 21088 11612 21100
rect 11664 21088 11670 21140
rect 15746 21088 15752 21140
rect 15804 21128 15810 21140
rect 18874 21128 18880 21140
rect 15804 21100 17540 21128
rect 18835 21100 18880 21128
rect 15804 21088 15810 21100
rect 7837 21063 7895 21069
rect 7837 21029 7849 21063
rect 7883 21029 7895 21063
rect 7837 21023 7895 21029
rect 7239 20964 7788 20992
rect 7239 20961 7251 20964
rect 7193 20955 7251 20961
rect 7377 20927 7435 20933
rect 7377 20893 7389 20927
rect 7423 20924 7435 20927
rect 7852 20924 7880 21023
rect 9398 21020 9404 21072
rect 9456 21060 9462 21072
rect 10413 21063 10471 21069
rect 10413 21060 10425 21063
rect 9456 21032 10425 21060
rect 9456 21020 9462 21032
rect 10413 21029 10425 21032
rect 10459 21029 10471 21063
rect 10413 21023 10471 21029
rect 8110 20952 8116 21004
rect 8168 20992 8174 21004
rect 8481 20995 8539 21001
rect 8481 20992 8493 20995
rect 8168 20964 8493 20992
rect 8168 20952 8174 20964
rect 8481 20961 8493 20964
rect 8527 20992 8539 20995
rect 9953 20995 10011 21001
rect 9953 20992 9965 20995
rect 8527 20964 9965 20992
rect 8527 20961 8539 20964
rect 8481 20955 8539 20961
rect 9953 20961 9965 20964
rect 9999 20961 10011 20995
rect 11514 20992 11520 21004
rect 9953 20955 10011 20961
rect 10980 20964 11520 20992
rect 7423 20896 7880 20924
rect 7423 20893 7435 20896
rect 7377 20887 7435 20893
rect 8202 20884 8208 20936
rect 8260 20924 8266 20936
rect 8297 20927 8355 20933
rect 8297 20924 8309 20927
rect 8260 20896 8309 20924
rect 8260 20884 8266 20896
rect 8297 20893 8309 20896
rect 8343 20893 8355 20927
rect 9766 20924 9772 20936
rect 9727 20896 9772 20924
rect 8297 20887 8355 20893
rect 9766 20884 9772 20896
rect 9824 20884 9830 20936
rect 10870 20924 10876 20936
rect 10831 20896 10876 20924
rect 10870 20884 10876 20896
rect 10928 20884 10934 20936
rect 10980 20933 11008 20964
rect 11514 20952 11520 20964
rect 11572 20952 11578 21004
rect 15013 20995 15071 21001
rect 15013 20961 15025 20995
rect 15059 20992 15071 20995
rect 15764 20992 15792 21088
rect 15841 21063 15899 21069
rect 15841 21029 15853 21063
rect 15887 21060 15899 21063
rect 16758 21060 16764 21072
rect 15887 21032 16764 21060
rect 15887 21029 15899 21032
rect 15841 21023 15899 21029
rect 16758 21020 16764 21032
rect 16816 21020 16822 21072
rect 16853 21063 16911 21069
rect 16853 21029 16865 21063
rect 16899 21029 16911 21063
rect 16853 21023 16911 21029
rect 16298 20992 16304 21004
rect 15059 20964 15792 20992
rect 16259 20964 16304 20992
rect 15059 20961 15071 20964
rect 15013 20955 15071 20961
rect 16298 20952 16304 20964
rect 16356 20952 16362 21004
rect 10965 20927 11023 20933
rect 10965 20893 10977 20927
rect 11011 20893 11023 20927
rect 10965 20887 11023 20893
rect 11149 20927 11207 20933
rect 11149 20893 11161 20927
rect 11195 20924 11207 20927
rect 11425 20927 11483 20933
rect 11425 20924 11437 20927
rect 11195 20896 11437 20924
rect 11195 20893 11207 20896
rect 11149 20887 11207 20893
rect 11425 20893 11437 20896
rect 11471 20893 11483 20927
rect 11425 20887 11483 20893
rect 11885 20927 11943 20933
rect 11885 20893 11897 20927
rect 11931 20924 11943 20927
rect 12434 20924 12440 20936
rect 11931 20896 12440 20924
rect 11931 20893 11943 20896
rect 11885 20887 11943 20893
rect 12434 20884 12440 20896
rect 12492 20924 12498 20936
rect 13538 20924 13544 20936
rect 12492 20896 13544 20924
rect 12492 20884 12498 20896
rect 13538 20884 13544 20896
rect 13596 20884 13602 20936
rect 15286 20924 15292 20936
rect 15247 20896 15292 20924
rect 15286 20884 15292 20896
rect 15344 20884 15350 20936
rect 15657 20927 15715 20933
rect 15657 20893 15669 20927
rect 15703 20893 15715 20927
rect 16868 20924 16896 21023
rect 17512 21001 17540 21100
rect 18874 21088 18880 21100
rect 18932 21088 18938 21140
rect 19705 21131 19763 21137
rect 19705 21097 19717 21131
rect 19751 21128 19763 21131
rect 20254 21128 20260 21140
rect 19751 21100 20260 21128
rect 19751 21097 19763 21100
rect 19705 21091 19763 21097
rect 20254 21088 20260 21100
rect 20312 21088 20318 21140
rect 24029 21131 24087 21137
rect 24029 21097 24041 21131
rect 24075 21128 24087 21131
rect 28074 21128 28080 21140
rect 24075 21100 28080 21128
rect 24075 21097 24087 21100
rect 24029 21091 24087 21097
rect 28074 21088 28080 21100
rect 28132 21088 28138 21140
rect 19981 21063 20039 21069
rect 19981 21029 19993 21063
rect 20027 21029 20039 21063
rect 19981 21023 20039 21029
rect 17497 20995 17555 21001
rect 17497 20961 17509 20995
rect 17543 20961 17555 20995
rect 17497 20955 17555 20961
rect 18233 20995 18291 21001
rect 18233 20961 18245 20995
rect 18279 20961 18291 20995
rect 18414 20992 18420 21004
rect 18375 20964 18420 20992
rect 18233 20955 18291 20961
rect 17313 20927 17371 20933
rect 17313 20924 17325 20927
rect 16868 20896 17325 20924
rect 15657 20887 15715 20893
rect 17313 20893 17325 20896
rect 17359 20893 17371 20927
rect 17313 20887 17371 20893
rect 9030 20856 9036 20868
rect 8220 20828 9036 20856
rect 8220 20797 8248 20828
rect 9030 20816 9036 20828
rect 9088 20856 9094 20868
rect 9861 20859 9919 20865
rect 9861 20856 9873 20859
rect 9088 20828 9873 20856
rect 9088 20816 9094 20828
rect 9861 20825 9873 20828
rect 9907 20856 9919 20859
rect 11238 20856 11244 20868
rect 9907 20828 11244 20856
rect 9907 20825 9919 20828
rect 9861 20819 9919 20825
rect 11238 20816 11244 20828
rect 11296 20816 11302 20868
rect 11330 20816 11336 20868
rect 11388 20856 11394 20868
rect 12130 20859 12188 20865
rect 12130 20856 12142 20859
rect 11388 20828 12142 20856
rect 11388 20816 11394 20828
rect 12130 20825 12142 20828
rect 12176 20825 12188 20859
rect 15672 20856 15700 20887
rect 17129 20859 17187 20865
rect 17129 20856 17141 20859
rect 15672 20828 17141 20856
rect 12130 20819 12188 20825
rect 17129 20825 17141 20828
rect 17175 20825 17187 20859
rect 18248 20856 18276 20955
rect 18414 20952 18420 20964
rect 18472 20952 18478 21004
rect 19334 20952 19340 21004
rect 19392 20992 19398 21004
rect 19610 20992 19616 21004
rect 19392 20964 19616 20992
rect 19392 20952 19398 20964
rect 19610 20952 19616 20964
rect 19668 20952 19674 21004
rect 19521 20927 19579 20933
rect 19521 20893 19533 20927
rect 19567 20924 19579 20927
rect 19996 20924 20024 21023
rect 20533 20995 20591 21001
rect 20533 20961 20545 20995
rect 20579 20961 20591 20995
rect 20533 20955 20591 20961
rect 19567 20896 20024 20924
rect 19567 20893 19579 20896
rect 19521 20887 19579 20893
rect 20548 20868 20576 20955
rect 21266 20884 21272 20936
rect 21324 20924 21330 20936
rect 22106 20927 22164 20933
rect 22106 20924 22118 20927
rect 21324 20896 22118 20924
rect 21324 20884 21330 20896
rect 22106 20893 22118 20896
rect 22152 20893 22164 20927
rect 22106 20887 22164 20893
rect 22373 20927 22431 20933
rect 22373 20893 22385 20927
rect 22419 20924 22431 20927
rect 22649 20927 22707 20933
rect 22649 20924 22661 20927
rect 22419 20896 22661 20924
rect 22419 20893 22431 20896
rect 22373 20887 22431 20893
rect 22649 20893 22661 20896
rect 22695 20924 22707 20927
rect 23198 20924 23204 20936
rect 22695 20896 23204 20924
rect 22695 20893 22707 20896
rect 22649 20887 22707 20893
rect 23198 20884 23204 20896
rect 23256 20884 23262 20936
rect 19886 20856 19892 20868
rect 18248 20828 19892 20856
rect 17129 20819 17187 20825
rect 19886 20816 19892 20828
rect 19944 20856 19950 20868
rect 20530 20856 20536 20868
rect 19944 20828 20536 20856
rect 19944 20816 19950 20828
rect 20530 20816 20536 20828
rect 20588 20816 20594 20868
rect 22462 20816 22468 20868
rect 22520 20856 22526 20868
rect 22894 20859 22952 20865
rect 22894 20856 22906 20859
rect 22520 20828 22906 20856
rect 22520 20816 22526 20828
rect 22894 20825 22906 20828
rect 22940 20825 22952 20859
rect 22894 20819 22952 20825
rect 8205 20791 8263 20797
rect 8205 20757 8217 20791
rect 8251 20757 8263 20791
rect 8205 20751 8263 20757
rect 9401 20791 9459 20797
rect 9401 20757 9413 20791
rect 9447 20788 9459 20791
rect 9490 20788 9496 20800
rect 9447 20760 9496 20788
rect 9447 20757 9459 20760
rect 9401 20751 9459 20757
rect 9490 20748 9496 20760
rect 9548 20748 9554 20800
rect 12802 20748 12808 20800
rect 12860 20788 12866 20800
rect 13265 20791 13323 20797
rect 13265 20788 13277 20791
rect 12860 20760 13277 20788
rect 12860 20748 12866 20760
rect 13265 20757 13277 20760
rect 13311 20757 13323 20791
rect 13265 20751 13323 20757
rect 13446 20748 13452 20800
rect 13504 20788 13510 20800
rect 14093 20791 14151 20797
rect 14093 20788 14105 20791
rect 13504 20760 14105 20788
rect 13504 20748 13510 20760
rect 14093 20757 14105 20760
rect 14139 20757 14151 20791
rect 14093 20751 14151 20757
rect 16114 20748 16120 20800
rect 16172 20788 16178 20800
rect 16393 20791 16451 20797
rect 16393 20788 16405 20791
rect 16172 20760 16405 20788
rect 16172 20748 16178 20760
rect 16393 20757 16405 20760
rect 16439 20757 16451 20791
rect 16393 20751 16451 20757
rect 16485 20791 16543 20797
rect 16485 20757 16497 20791
rect 16531 20788 16543 20791
rect 17865 20791 17923 20797
rect 17865 20788 17877 20791
rect 16531 20760 17877 20788
rect 16531 20757 16543 20760
rect 16485 20751 16543 20757
rect 17865 20757 17877 20760
rect 17911 20788 17923 20791
rect 18509 20791 18567 20797
rect 18509 20788 18521 20791
rect 17911 20760 18521 20788
rect 17911 20757 17923 20760
rect 17865 20751 17923 20757
rect 18509 20757 18521 20760
rect 18555 20788 18567 20791
rect 19242 20788 19248 20800
rect 18555 20760 19248 20788
rect 18555 20757 18567 20760
rect 18509 20751 18567 20757
rect 19242 20748 19248 20760
rect 19300 20748 19306 20800
rect 20254 20748 20260 20800
rect 20312 20788 20318 20800
rect 20349 20791 20407 20797
rect 20349 20788 20361 20791
rect 20312 20760 20361 20788
rect 20312 20748 20318 20760
rect 20349 20757 20361 20760
rect 20395 20757 20407 20791
rect 20349 20751 20407 20757
rect 20438 20748 20444 20800
rect 20496 20788 20502 20800
rect 20993 20791 21051 20797
rect 20993 20788 21005 20791
rect 20496 20760 21005 20788
rect 20496 20748 20502 20760
rect 20993 20757 21005 20760
rect 21039 20757 21051 20791
rect 20993 20751 21051 20757
rect 1104 20698 28888 20720
rect 1104 20646 10214 20698
rect 10266 20646 10278 20698
rect 10330 20646 10342 20698
rect 10394 20646 10406 20698
rect 10458 20646 10470 20698
rect 10522 20646 19478 20698
rect 19530 20646 19542 20698
rect 19594 20646 19606 20698
rect 19658 20646 19670 20698
rect 19722 20646 19734 20698
rect 19786 20646 28888 20698
rect 1104 20624 28888 20646
rect 9674 20584 9680 20596
rect 9635 20556 9680 20584
rect 9674 20544 9680 20556
rect 9732 20544 9738 20596
rect 11146 20584 11152 20596
rect 11107 20556 11152 20584
rect 11146 20544 11152 20556
rect 11204 20544 11210 20596
rect 11238 20544 11244 20596
rect 11296 20584 11302 20596
rect 12253 20587 12311 20593
rect 12253 20584 12265 20587
rect 11296 20556 12265 20584
rect 11296 20544 11302 20556
rect 12253 20553 12265 20556
rect 12299 20553 12311 20587
rect 12253 20547 12311 20553
rect 15013 20587 15071 20593
rect 15013 20553 15025 20587
rect 15059 20584 15071 20587
rect 15470 20584 15476 20596
rect 15059 20556 15476 20584
rect 15059 20553 15071 20556
rect 15013 20547 15071 20553
rect 15470 20544 15476 20556
rect 15528 20584 15534 20596
rect 15528 20556 17264 20584
rect 15528 20544 15534 20556
rect 8941 20519 8999 20525
rect 8941 20485 8953 20519
rect 8987 20516 8999 20519
rect 10134 20516 10140 20528
rect 8987 20488 10140 20516
rect 8987 20485 8999 20488
rect 8941 20479 8999 20485
rect 10134 20476 10140 20488
rect 10192 20516 10198 20528
rect 13265 20519 13323 20525
rect 13265 20516 13277 20519
rect 10192 20488 13277 20516
rect 10192 20476 10198 20488
rect 13265 20485 13277 20488
rect 13311 20485 13323 20519
rect 13265 20479 13323 20485
rect 15841 20519 15899 20525
rect 15841 20485 15853 20519
rect 15887 20516 15899 20519
rect 16298 20516 16304 20528
rect 15887 20488 16304 20516
rect 15887 20485 15899 20488
rect 15841 20479 15899 20485
rect 7098 20457 7104 20460
rect 7092 20411 7104 20457
rect 7156 20448 7162 20460
rect 9490 20448 9496 20460
rect 7156 20420 7192 20448
rect 9451 20420 9496 20448
rect 7098 20408 7104 20411
rect 7156 20408 7162 20420
rect 9490 20408 9496 20420
rect 9548 20408 9554 20460
rect 10042 20408 10048 20460
rect 10100 20448 10106 20460
rect 10321 20451 10379 20457
rect 10321 20448 10333 20451
rect 10100 20420 10333 20448
rect 10100 20408 10106 20420
rect 10321 20417 10333 20420
rect 10367 20417 10379 20451
rect 10870 20448 10876 20460
rect 10831 20420 10876 20448
rect 10321 20411 10379 20417
rect 10870 20408 10876 20420
rect 10928 20408 10934 20460
rect 10965 20451 11023 20457
rect 10965 20417 10977 20451
rect 11011 20448 11023 20451
rect 12161 20451 12219 20457
rect 11011 20420 11836 20448
rect 11011 20417 11023 20420
rect 10965 20411 11023 20417
rect 6822 20380 6828 20392
rect 6783 20352 6828 20380
rect 6822 20340 6828 20352
rect 6880 20340 6886 20392
rect 9309 20383 9367 20389
rect 9309 20349 9321 20383
rect 9355 20380 9367 20383
rect 9398 20380 9404 20392
rect 9355 20352 9404 20380
rect 9355 20349 9367 20352
rect 9309 20343 9367 20349
rect 9398 20340 9404 20352
rect 9456 20340 9462 20392
rect 10137 20383 10195 20389
rect 10137 20349 10149 20383
rect 10183 20380 10195 20383
rect 10888 20380 10916 20408
rect 10183 20352 10916 20380
rect 10183 20349 10195 20352
rect 10137 20343 10195 20349
rect 11808 20321 11836 20420
rect 12161 20417 12173 20451
rect 12207 20448 12219 20451
rect 12802 20448 12808 20460
rect 12207 20420 12808 20448
rect 12207 20417 12219 20420
rect 12161 20411 12219 20417
rect 12802 20408 12808 20420
rect 12860 20408 12866 20460
rect 13630 20408 13636 20460
rect 13688 20448 13694 20460
rect 13725 20451 13783 20457
rect 13725 20448 13737 20451
rect 13688 20420 13737 20448
rect 13688 20408 13694 20420
rect 13725 20417 13737 20420
rect 13771 20417 13783 20451
rect 14274 20448 14280 20460
rect 14235 20420 14280 20448
rect 13725 20411 13783 20417
rect 14274 20408 14280 20420
rect 14332 20448 14338 20460
rect 14921 20451 14979 20457
rect 14921 20448 14933 20451
rect 14332 20420 14933 20448
rect 14332 20408 14338 20420
rect 14921 20417 14933 20420
rect 14967 20417 14979 20451
rect 14921 20411 14979 20417
rect 15562 20408 15568 20460
rect 15620 20448 15626 20460
rect 15657 20451 15715 20457
rect 15657 20448 15669 20451
rect 15620 20420 15669 20448
rect 15620 20408 15626 20420
rect 15657 20417 15669 20420
rect 15703 20417 15715 20451
rect 15657 20411 15715 20417
rect 12342 20380 12348 20392
rect 12303 20352 12348 20380
rect 12342 20340 12348 20352
rect 12400 20340 12406 20392
rect 15197 20383 15255 20389
rect 15197 20349 15209 20383
rect 15243 20380 15255 20383
rect 15856 20380 15884 20479
rect 16298 20476 16304 20488
rect 16356 20476 16362 20528
rect 17126 20516 17132 20528
rect 16684 20488 17132 20516
rect 16684 20457 16712 20488
rect 17126 20476 17132 20488
rect 17184 20476 17190 20528
rect 17236 20516 17264 20556
rect 18322 20544 18328 20596
rect 18380 20584 18386 20596
rect 18509 20587 18567 20593
rect 18509 20584 18521 20587
rect 18380 20556 18521 20584
rect 18380 20544 18386 20556
rect 18509 20553 18521 20556
rect 18555 20553 18567 20587
rect 18509 20547 18567 20553
rect 19334 20544 19340 20596
rect 19392 20584 19398 20596
rect 19613 20587 19671 20593
rect 19613 20584 19625 20587
rect 19392 20556 19625 20584
rect 19392 20544 19398 20556
rect 19613 20553 19625 20556
rect 19659 20553 19671 20587
rect 19613 20547 19671 20553
rect 19889 20587 19947 20593
rect 19889 20553 19901 20587
rect 19935 20584 19947 20587
rect 20162 20584 20168 20596
rect 19935 20556 20168 20584
rect 19935 20553 19947 20556
rect 19889 20547 19947 20553
rect 20162 20544 20168 20556
rect 20220 20544 20226 20596
rect 21085 20587 21143 20593
rect 21085 20553 21097 20587
rect 21131 20584 21143 20587
rect 21131 20556 22094 20584
rect 21131 20553 21143 20556
rect 21085 20547 21143 20553
rect 18877 20519 18935 20525
rect 18877 20516 18889 20519
rect 17236 20488 18889 20516
rect 18877 20485 18889 20488
rect 18923 20485 18935 20519
rect 20438 20516 20444 20528
rect 18877 20479 18935 20485
rect 19076 20488 20444 20516
rect 16669 20451 16727 20457
rect 16669 20417 16681 20451
rect 16715 20417 16727 20451
rect 16669 20411 16727 20417
rect 16758 20408 16764 20460
rect 16816 20448 16822 20460
rect 16925 20451 16983 20457
rect 16925 20448 16937 20451
rect 16816 20420 16937 20448
rect 16816 20408 16822 20420
rect 16925 20417 16937 20420
rect 16971 20417 16983 20451
rect 16925 20411 16983 20417
rect 18688 20451 18746 20457
rect 18688 20417 18700 20451
rect 18734 20417 18746 20451
rect 18688 20411 18746 20417
rect 15243 20352 15884 20380
rect 18708 20380 18736 20411
rect 18782 20408 18788 20460
rect 18840 20448 18846 20460
rect 19076 20457 19104 20488
rect 20438 20476 20444 20488
rect 20496 20476 20502 20528
rect 22066 20516 22094 20556
rect 22934 20519 22992 20525
rect 22934 20516 22946 20519
rect 22066 20488 22946 20516
rect 22934 20485 22946 20488
rect 22980 20485 22992 20519
rect 22934 20479 22992 20485
rect 19060 20451 19118 20457
rect 18840 20420 18885 20448
rect 18840 20408 18846 20420
rect 19060 20417 19072 20451
rect 19106 20417 19118 20451
rect 19060 20411 19118 20417
rect 19150 20408 19156 20460
rect 19208 20448 19214 20460
rect 19429 20451 19487 20457
rect 19208 20420 19253 20448
rect 19208 20408 19214 20420
rect 19429 20417 19441 20451
rect 19475 20448 19487 20451
rect 19978 20448 19984 20460
rect 19475 20420 19984 20448
rect 19475 20417 19487 20420
rect 19429 20411 19487 20417
rect 19978 20408 19984 20420
rect 20036 20408 20042 20460
rect 20162 20408 20168 20460
rect 20220 20448 20226 20460
rect 20257 20451 20315 20457
rect 20257 20448 20269 20451
rect 20220 20420 20269 20448
rect 20220 20408 20226 20420
rect 20257 20417 20269 20420
rect 20303 20417 20315 20451
rect 20898 20448 20904 20460
rect 20859 20420 20904 20448
rect 20257 20411 20315 20417
rect 20898 20408 20904 20420
rect 20956 20408 20962 20460
rect 20349 20383 20407 20389
rect 20349 20380 20361 20383
rect 18708 20352 20361 20380
rect 15243 20349 15255 20352
rect 15197 20343 15255 20349
rect 20349 20349 20361 20352
rect 20395 20349 20407 20383
rect 20530 20380 20536 20392
rect 20491 20352 20536 20380
rect 20349 20343 20407 20349
rect 11793 20315 11851 20321
rect 11793 20281 11805 20315
rect 11839 20281 11851 20315
rect 11793 20275 11851 20281
rect 13449 20315 13507 20321
rect 13449 20281 13461 20315
rect 13495 20312 13507 20315
rect 13538 20312 13544 20324
rect 13495 20284 13544 20312
rect 13495 20281 13507 20284
rect 13449 20275 13507 20281
rect 13538 20272 13544 20284
rect 13596 20272 13602 20324
rect 20364 20312 20392 20343
rect 20530 20340 20536 20352
rect 20588 20340 20594 20392
rect 23198 20380 23204 20392
rect 23159 20352 23204 20380
rect 23198 20340 23204 20352
rect 23256 20340 23262 20392
rect 21821 20315 21879 20321
rect 21821 20312 21833 20315
rect 20364 20284 21833 20312
rect 21821 20281 21833 20284
rect 21867 20281 21879 20315
rect 21821 20275 21879 20281
rect 8202 20244 8208 20256
rect 8163 20216 8208 20244
rect 8202 20204 8208 20216
rect 8260 20204 8266 20256
rect 8849 20247 8907 20253
rect 8849 20213 8861 20247
rect 8895 20244 8907 20247
rect 9122 20244 9128 20256
rect 8895 20216 9128 20244
rect 8895 20213 8907 20216
rect 8849 20207 8907 20213
rect 9122 20204 9128 20216
rect 9180 20204 9186 20256
rect 10505 20247 10563 20253
rect 10505 20213 10517 20247
rect 10551 20244 10563 20247
rect 11698 20244 11704 20256
rect 10551 20216 11704 20244
rect 10551 20213 10563 20216
rect 10505 20207 10563 20213
rect 11698 20204 11704 20216
rect 11756 20204 11762 20256
rect 13906 20244 13912 20256
rect 13867 20216 13912 20244
rect 13906 20204 13912 20216
rect 13964 20204 13970 20256
rect 14550 20244 14556 20256
rect 14511 20216 14556 20244
rect 14550 20204 14556 20216
rect 14608 20204 14614 20256
rect 16114 20204 16120 20256
rect 16172 20244 16178 20256
rect 18049 20247 18107 20253
rect 18049 20244 18061 20247
rect 16172 20216 18061 20244
rect 16172 20204 16178 20216
rect 18049 20213 18061 20216
rect 18095 20244 18107 20247
rect 18414 20244 18420 20256
rect 18095 20216 18420 20244
rect 18095 20213 18107 20216
rect 18049 20207 18107 20213
rect 18414 20204 18420 20216
rect 18472 20204 18478 20256
rect 1104 20154 28888 20176
rect 1104 20102 5582 20154
rect 5634 20102 5646 20154
rect 5698 20102 5710 20154
rect 5762 20102 5774 20154
rect 5826 20102 5838 20154
rect 5890 20102 14846 20154
rect 14898 20102 14910 20154
rect 14962 20102 14974 20154
rect 15026 20102 15038 20154
rect 15090 20102 15102 20154
rect 15154 20102 24110 20154
rect 24162 20102 24174 20154
rect 24226 20102 24238 20154
rect 24290 20102 24302 20154
rect 24354 20102 24366 20154
rect 24418 20102 28888 20154
rect 1104 20080 28888 20102
rect 6917 20043 6975 20049
rect 6917 20009 6929 20043
rect 6963 20040 6975 20043
rect 7098 20040 7104 20052
rect 6963 20012 7104 20040
rect 6963 20009 6975 20012
rect 6917 20003 6975 20009
rect 7098 20000 7104 20012
rect 7156 20000 7162 20052
rect 12342 20000 12348 20052
rect 12400 20040 12406 20052
rect 15470 20040 15476 20052
rect 12400 20012 15332 20040
rect 15431 20012 15476 20040
rect 12400 20000 12406 20012
rect 7837 19975 7895 19981
rect 7837 19941 7849 19975
rect 7883 19941 7895 19975
rect 7837 19935 7895 19941
rect 7852 19904 7880 19935
rect 7392 19876 7880 19904
rect 1394 19836 1400 19848
rect 1355 19808 1400 19836
rect 1394 19796 1400 19808
rect 1452 19796 1458 19848
rect 7392 19845 7420 19876
rect 8110 19864 8116 19916
rect 8168 19904 8174 19916
rect 8389 19907 8447 19913
rect 8389 19904 8401 19907
rect 8168 19876 8401 19904
rect 8168 19864 8174 19876
rect 8389 19873 8401 19876
rect 8435 19873 8447 19907
rect 8389 19867 8447 19873
rect 13538 19864 13544 19916
rect 13596 19904 13602 19916
rect 14093 19907 14151 19913
rect 14093 19904 14105 19907
rect 13596 19876 14105 19904
rect 13596 19864 13602 19876
rect 14093 19873 14105 19876
rect 14139 19873 14151 19907
rect 15304 19904 15332 20012
rect 15470 20000 15476 20012
rect 15528 20000 15534 20052
rect 16206 20000 16212 20052
rect 16264 20040 16270 20052
rect 17129 20043 17187 20049
rect 17129 20040 17141 20043
rect 16264 20012 17141 20040
rect 16264 20000 16270 20012
rect 17129 20009 17141 20012
rect 17175 20009 17187 20043
rect 17129 20003 17187 20009
rect 18601 20043 18659 20049
rect 18601 20009 18613 20043
rect 18647 20040 18659 20043
rect 19150 20040 19156 20052
rect 18647 20012 19156 20040
rect 18647 20009 18659 20012
rect 18601 20003 18659 20009
rect 19150 20000 19156 20012
rect 19208 20000 19214 20052
rect 19242 20000 19248 20052
rect 19300 20040 19306 20052
rect 19337 20043 19395 20049
rect 19337 20040 19349 20043
rect 19300 20012 19349 20040
rect 19300 20000 19306 20012
rect 19337 20009 19349 20012
rect 19383 20040 19395 20043
rect 22738 20040 22744 20052
rect 19383 20012 22744 20040
rect 19383 20009 19395 20012
rect 19337 20003 19395 20009
rect 22738 20000 22744 20012
rect 22796 20000 22802 20052
rect 20070 19932 20076 19984
rect 20128 19972 20134 19984
rect 21453 19975 21511 19981
rect 21453 19972 21465 19975
rect 20128 19944 21465 19972
rect 20128 19932 20134 19944
rect 21453 19941 21465 19944
rect 21499 19972 21511 19975
rect 21499 19944 22232 19972
rect 21499 19941 21511 19944
rect 21453 19935 21511 19941
rect 19886 19904 19892 19916
rect 15304 19876 17080 19904
rect 14093 19867 14151 19873
rect 1673 19839 1731 19845
rect 1673 19805 1685 19839
rect 1719 19805 1731 19839
rect 1673 19799 1731 19805
rect 6733 19839 6791 19845
rect 6733 19805 6745 19839
rect 6779 19836 6791 19839
rect 7193 19839 7251 19845
rect 7193 19836 7205 19839
rect 6779 19808 7205 19836
rect 6779 19805 6791 19808
rect 6733 19799 6791 19805
rect 7193 19805 7205 19808
rect 7239 19805 7251 19839
rect 7193 19799 7251 19805
rect 7377 19839 7435 19845
rect 7377 19805 7389 19839
rect 7423 19805 7435 19839
rect 7377 19799 7435 19805
rect 7561 19839 7619 19845
rect 7561 19805 7573 19839
rect 7607 19836 7619 19839
rect 8294 19836 8300 19848
rect 7607 19808 8300 19836
rect 7607 19805 7619 19808
rect 7561 19799 7619 19805
rect 1688 19768 1716 19799
rect 8294 19796 8300 19808
rect 8352 19796 8358 19848
rect 9030 19836 9036 19848
rect 8991 19808 9036 19836
rect 9030 19796 9036 19808
rect 9088 19796 9094 19848
rect 9122 19796 9128 19848
rect 9180 19836 9186 19848
rect 10965 19839 11023 19845
rect 10965 19836 10977 19839
rect 9180 19808 10977 19836
rect 9180 19796 9186 19808
rect 10965 19805 10977 19808
rect 11011 19805 11023 19839
rect 10965 19799 11023 19805
rect 13078 19796 13084 19848
rect 13136 19836 13142 19848
rect 13449 19839 13507 19845
rect 13449 19836 13461 19839
rect 13136 19808 13461 19836
rect 13136 19796 13142 19808
rect 13449 19805 13461 19808
rect 13495 19805 13507 19839
rect 13449 19799 13507 19805
rect 13725 19839 13783 19845
rect 13725 19805 13737 19839
rect 13771 19805 13783 19839
rect 13725 19799 13783 19805
rect 7742 19768 7748 19780
rect 1688 19740 7748 19768
rect 7742 19728 7748 19740
rect 7800 19728 7806 19780
rect 9306 19777 9312 19780
rect 9300 19731 9312 19777
rect 9364 19768 9370 19780
rect 11232 19771 11290 19777
rect 9364 19740 9400 19768
rect 9306 19728 9312 19731
rect 9364 19728 9370 19740
rect 11232 19737 11244 19771
rect 11278 19768 11290 19771
rect 11514 19768 11520 19780
rect 11278 19740 11520 19768
rect 11278 19737 11290 19740
rect 11232 19731 11290 19737
rect 11514 19728 11520 19740
rect 11572 19728 11578 19780
rect 13740 19768 13768 19799
rect 13906 19796 13912 19848
rect 13964 19836 13970 19848
rect 14349 19839 14407 19845
rect 14349 19836 14361 19839
rect 13964 19808 14361 19836
rect 13964 19796 13970 19808
rect 14349 19805 14361 19808
rect 14395 19805 14407 19839
rect 14349 19799 14407 19805
rect 15933 19839 15991 19845
rect 15933 19805 15945 19839
rect 15979 19805 15991 19839
rect 16114 19836 16120 19848
rect 16075 19808 16120 19836
rect 15933 19799 15991 19805
rect 15286 19768 15292 19780
rect 13740 19740 15292 19768
rect 15286 19728 15292 19740
rect 15344 19728 15350 19780
rect 15948 19768 15976 19799
rect 16114 19796 16120 19808
rect 16172 19796 16178 19848
rect 16209 19839 16267 19845
rect 16209 19805 16221 19839
rect 16255 19836 16267 19839
rect 16574 19836 16580 19848
rect 16255 19808 16580 19836
rect 16255 19805 16267 19808
rect 16209 19799 16267 19805
rect 16574 19796 16580 19808
rect 16632 19796 16638 19848
rect 17052 19845 17080 19876
rect 18156 19876 19892 19904
rect 17037 19839 17095 19845
rect 17037 19805 17049 19839
rect 17083 19836 17095 19839
rect 17678 19836 17684 19848
rect 17083 19808 17684 19836
rect 17083 19805 17095 19808
rect 17037 19799 17095 19805
rect 17678 19796 17684 19808
rect 17736 19796 17742 19848
rect 17954 19836 17960 19848
rect 17915 19808 17960 19836
rect 17954 19796 17960 19808
rect 18012 19796 18018 19848
rect 18156 19845 18184 19876
rect 19886 19864 19892 19876
rect 19944 19864 19950 19916
rect 20254 19864 20260 19916
rect 20312 19904 20318 19916
rect 22005 19907 22063 19913
rect 22005 19904 22017 19907
rect 20312 19876 22017 19904
rect 20312 19864 20318 19876
rect 22005 19873 22017 19876
rect 22051 19904 22063 19907
rect 22094 19904 22100 19916
rect 22051 19876 22100 19904
rect 22051 19873 22063 19876
rect 22005 19867 22063 19873
rect 22094 19864 22100 19876
rect 22152 19864 22158 19916
rect 22204 19904 22232 19944
rect 22204 19876 22508 19904
rect 18105 19839 18184 19845
rect 18105 19805 18117 19839
rect 18151 19808 18184 19839
rect 18322 19836 18328 19848
rect 18283 19808 18328 19836
rect 18151 19805 18163 19808
rect 18105 19799 18163 19805
rect 18322 19796 18328 19808
rect 18380 19796 18386 19848
rect 18414 19796 18420 19848
rect 18472 19845 18478 19848
rect 18472 19836 18480 19845
rect 18472 19808 18517 19836
rect 18472 19799 18480 19808
rect 18472 19796 18478 19799
rect 20622 19796 20628 19848
rect 20680 19836 20686 19848
rect 22373 19839 22431 19845
rect 22373 19836 22385 19839
rect 20680 19808 22385 19836
rect 20680 19796 20686 19808
rect 22373 19805 22385 19808
rect 22419 19805 22431 19839
rect 22480 19836 22508 19876
rect 24210 19836 24216 19848
rect 22480 19808 24216 19836
rect 22373 19799 22431 19805
rect 24210 19796 24216 19808
rect 24268 19796 24274 19848
rect 16022 19768 16028 19780
rect 15580 19740 15884 19768
rect 15948 19740 16028 19768
rect 8202 19700 8208 19712
rect 8163 19672 8208 19700
rect 8202 19660 8208 19672
rect 8260 19660 8266 19712
rect 8297 19703 8355 19709
rect 8297 19669 8309 19703
rect 8343 19700 8355 19703
rect 9674 19700 9680 19712
rect 8343 19672 9680 19700
rect 8343 19669 8355 19672
rect 8297 19663 8355 19669
rect 9674 19660 9680 19672
rect 9732 19700 9738 19712
rect 10413 19703 10471 19709
rect 10413 19700 10425 19703
rect 9732 19672 10425 19700
rect 9732 19660 9738 19672
rect 10413 19669 10425 19672
rect 10459 19669 10471 19703
rect 10413 19663 10471 19669
rect 12250 19660 12256 19712
rect 12308 19700 12314 19712
rect 12345 19703 12403 19709
rect 12345 19700 12357 19703
rect 12308 19672 12357 19700
rect 12308 19660 12314 19672
rect 12345 19669 12357 19672
rect 12391 19669 12403 19703
rect 12345 19663 12403 19669
rect 14274 19660 14280 19712
rect 14332 19700 14338 19712
rect 15580 19700 15608 19740
rect 15746 19700 15752 19712
rect 14332 19672 15608 19700
rect 15707 19672 15752 19700
rect 14332 19660 14338 19672
rect 15746 19660 15752 19672
rect 15804 19660 15810 19712
rect 15856 19700 15884 19740
rect 16022 19728 16028 19740
rect 16080 19728 16086 19780
rect 18230 19768 18236 19780
rect 17328 19740 17632 19768
rect 18191 19740 18236 19768
rect 17328 19700 17356 19740
rect 15856 19672 17356 19700
rect 17402 19660 17408 19712
rect 17460 19700 17466 19712
rect 17497 19703 17555 19709
rect 17497 19700 17509 19703
rect 17460 19672 17509 19700
rect 17460 19660 17466 19672
rect 17497 19669 17509 19672
rect 17543 19669 17555 19703
rect 17604 19700 17632 19740
rect 18230 19728 18236 19740
rect 18288 19728 18294 19780
rect 20073 19771 20131 19777
rect 20073 19768 20085 19771
rect 19720 19740 20085 19768
rect 19720 19700 19748 19740
rect 20073 19737 20085 19740
rect 20119 19768 20131 19771
rect 20254 19768 20260 19780
rect 20119 19740 20260 19768
rect 20119 19737 20131 19740
rect 20073 19731 20131 19737
rect 20254 19728 20260 19740
rect 20312 19728 20318 19780
rect 21637 19771 21695 19777
rect 21637 19737 21649 19771
rect 21683 19737 21695 19771
rect 21637 19731 21695 19737
rect 17604 19672 19748 19700
rect 19797 19703 19855 19709
rect 17497 19663 17555 19669
rect 19797 19669 19809 19703
rect 19843 19700 19855 19703
rect 20162 19700 20168 19712
rect 19843 19672 20168 19700
rect 19843 19669 19855 19672
rect 19797 19663 19855 19669
rect 20162 19660 20168 19672
rect 20220 19700 20226 19712
rect 20530 19700 20536 19712
rect 20220 19672 20536 19700
rect 20220 19660 20226 19672
rect 20530 19660 20536 19672
rect 20588 19660 20594 19712
rect 21082 19700 21088 19712
rect 21043 19672 21088 19700
rect 21082 19660 21088 19672
rect 21140 19700 21146 19712
rect 21652 19700 21680 19731
rect 21726 19728 21732 19780
rect 21784 19768 21790 19780
rect 22646 19777 22652 19780
rect 21784 19740 22600 19768
rect 21784 19728 21790 19740
rect 21140 19672 21680 19700
rect 22572 19700 22600 19740
rect 22640 19731 22652 19777
rect 22704 19768 22710 19780
rect 22704 19740 22740 19768
rect 22646 19728 22652 19731
rect 22704 19728 22710 19740
rect 23014 19700 23020 19712
rect 22572 19672 23020 19700
rect 21140 19660 21146 19672
rect 23014 19660 23020 19672
rect 23072 19700 23078 19712
rect 23753 19703 23811 19709
rect 23753 19700 23765 19703
rect 23072 19672 23765 19700
rect 23072 19660 23078 19672
rect 23753 19669 23765 19672
rect 23799 19669 23811 19703
rect 23753 19663 23811 19669
rect 1104 19610 28888 19632
rect 1104 19558 10214 19610
rect 10266 19558 10278 19610
rect 10330 19558 10342 19610
rect 10394 19558 10406 19610
rect 10458 19558 10470 19610
rect 10522 19558 19478 19610
rect 19530 19558 19542 19610
rect 19594 19558 19606 19610
rect 19658 19558 19670 19610
rect 19722 19558 19734 19610
rect 19786 19558 28888 19610
rect 1104 19536 28888 19558
rect 1394 19496 1400 19508
rect 1355 19468 1400 19496
rect 1394 19456 1400 19468
rect 1452 19456 1458 19508
rect 6825 19499 6883 19505
rect 6825 19465 6837 19499
rect 6871 19496 6883 19499
rect 6914 19496 6920 19508
rect 6871 19468 6920 19496
rect 6871 19465 6883 19468
rect 6825 19459 6883 19465
rect 6914 19456 6920 19468
rect 6972 19456 6978 19508
rect 9306 19496 9312 19508
rect 9267 19468 9312 19496
rect 9306 19456 9312 19468
rect 9364 19456 9370 19508
rect 10042 19456 10048 19508
rect 10100 19496 10106 19508
rect 10413 19499 10471 19505
rect 10413 19496 10425 19499
rect 10100 19468 10425 19496
rect 10100 19456 10106 19468
rect 10413 19465 10425 19468
rect 10459 19465 10471 19499
rect 11514 19496 11520 19508
rect 11475 19468 11520 19496
rect 10413 19459 10471 19465
rect 11514 19456 11520 19468
rect 11572 19456 11578 19508
rect 13630 19496 13636 19508
rect 13591 19468 13636 19496
rect 13630 19456 13636 19468
rect 13688 19456 13694 19508
rect 15470 19496 15476 19508
rect 15431 19468 15476 19496
rect 15470 19456 15476 19468
rect 15528 19456 15534 19508
rect 16206 19496 16212 19508
rect 16167 19468 16212 19496
rect 16206 19456 16212 19468
rect 16264 19496 16270 19508
rect 16264 19468 16988 19496
rect 16264 19456 16270 19468
rect 8202 19388 8208 19440
rect 8260 19428 8266 19440
rect 10781 19431 10839 19437
rect 8260 19400 9628 19428
rect 8260 19388 8266 19400
rect 7006 19360 7012 19372
rect 6967 19332 7012 19360
rect 7006 19320 7012 19332
rect 7064 19320 7070 19372
rect 8846 19360 8852 19372
rect 8807 19332 8852 19360
rect 8846 19320 8852 19332
rect 8904 19320 8910 19372
rect 9033 19363 9091 19369
rect 9033 19329 9045 19363
rect 9079 19360 9091 19363
rect 9493 19363 9551 19369
rect 9493 19360 9505 19363
rect 9079 19332 9505 19360
rect 9079 19329 9091 19332
rect 9033 19323 9091 19329
rect 9493 19329 9505 19332
rect 9539 19329 9551 19363
rect 9600 19360 9628 19400
rect 10781 19397 10793 19431
rect 10827 19428 10839 19431
rect 12250 19428 12256 19440
rect 10827 19400 12256 19428
rect 10827 19397 10839 19400
rect 10781 19391 10839 19397
rect 12250 19388 12256 19400
rect 12308 19388 12314 19440
rect 16960 19428 16988 19468
rect 17034 19456 17040 19508
rect 17092 19496 17098 19508
rect 18782 19496 18788 19508
rect 17092 19468 17137 19496
rect 17420 19468 18788 19496
rect 17092 19456 17098 19468
rect 17420 19428 17448 19468
rect 18782 19456 18788 19468
rect 18840 19496 18846 19508
rect 18877 19499 18935 19505
rect 18877 19496 18889 19499
rect 18840 19468 18889 19496
rect 18840 19456 18846 19468
rect 18877 19465 18889 19468
rect 18923 19465 18935 19499
rect 20438 19496 20444 19508
rect 18877 19459 18935 19465
rect 19628 19468 20444 19496
rect 19628 19440 19656 19468
rect 20438 19456 20444 19468
rect 20496 19456 20502 19508
rect 22557 19499 22615 19505
rect 22066 19468 22324 19496
rect 19334 19428 19340 19440
rect 15304 19400 16896 19428
rect 16960 19400 17448 19428
rect 17512 19400 19340 19428
rect 10873 19363 10931 19369
rect 10873 19360 10885 19363
rect 9600 19332 10885 19360
rect 9493 19323 9551 19329
rect 10873 19329 10885 19332
rect 10919 19329 10931 19363
rect 11698 19360 11704 19372
rect 11659 19332 11704 19360
rect 10873 19323 10931 19329
rect 11698 19320 11704 19332
rect 11756 19320 11762 19372
rect 12437 19363 12495 19369
rect 12437 19329 12449 19363
rect 12483 19360 12495 19363
rect 12526 19360 12532 19372
rect 12483 19332 12532 19360
rect 12483 19329 12495 19332
rect 12437 19323 12495 19329
rect 12526 19320 12532 19332
rect 12584 19320 12590 19372
rect 13449 19363 13507 19369
rect 13449 19329 13461 19363
rect 13495 19360 13507 19363
rect 14550 19360 14556 19372
rect 13495 19332 14556 19360
rect 13495 19329 13507 19332
rect 13449 19323 13507 19329
rect 14550 19320 14556 19332
rect 14608 19320 14614 19372
rect 15304 19369 15332 19400
rect 16040 19372 16068 19400
rect 15289 19363 15347 19369
rect 15289 19329 15301 19363
rect 15335 19329 15347 19363
rect 15289 19323 15347 19329
rect 15565 19363 15623 19369
rect 15565 19329 15577 19363
rect 15611 19329 15623 19363
rect 16022 19360 16028 19372
rect 15983 19332 16028 19360
rect 15565 19323 15623 19329
rect 7745 19295 7803 19301
rect 7745 19261 7757 19295
rect 7791 19292 7803 19295
rect 8294 19292 8300 19304
rect 7791 19264 8300 19292
rect 7791 19261 7803 19264
rect 7745 19255 7803 19261
rect 8294 19252 8300 19264
rect 8352 19292 8358 19304
rect 8665 19295 8723 19301
rect 8665 19292 8677 19295
rect 8352 19264 8677 19292
rect 8352 19252 8358 19264
rect 8665 19261 8677 19264
rect 8711 19292 8723 19295
rect 9398 19292 9404 19304
rect 8711 19264 9404 19292
rect 8711 19261 8723 19264
rect 8665 19255 8723 19261
rect 9398 19252 9404 19264
rect 9456 19292 9462 19304
rect 9861 19295 9919 19301
rect 9861 19292 9873 19295
rect 9456 19264 9873 19292
rect 9456 19252 9462 19264
rect 9861 19261 9873 19264
rect 9907 19292 9919 19295
rect 10962 19292 10968 19304
rect 9907 19264 9996 19292
rect 10923 19264 10968 19292
rect 9907 19261 9919 19264
rect 9861 19255 9919 19261
rect 9968 19224 9996 19264
rect 10962 19252 10968 19264
rect 11020 19252 11026 19304
rect 11238 19252 11244 19304
rect 11296 19292 11302 19304
rect 12161 19295 12219 19301
rect 12161 19292 12173 19295
rect 11296 19264 12173 19292
rect 11296 19252 11302 19264
rect 12161 19261 12173 19264
rect 12207 19261 12219 19295
rect 12161 19255 12219 19261
rect 13078 19252 13084 19304
rect 13136 19292 13142 19304
rect 13265 19295 13323 19301
rect 13265 19292 13277 19295
rect 13136 19264 13277 19292
rect 13136 19252 13142 19264
rect 13265 19261 13277 19264
rect 13311 19261 13323 19295
rect 13265 19255 13323 19261
rect 14642 19252 14648 19304
rect 14700 19292 14706 19304
rect 14737 19295 14795 19301
rect 14737 19292 14749 19295
rect 14700 19264 14749 19292
rect 14700 19252 14706 19264
rect 14737 19261 14749 19264
rect 14783 19261 14795 19295
rect 15580 19292 15608 19323
rect 16022 19320 16028 19332
rect 16080 19320 16086 19372
rect 16301 19363 16359 19369
rect 16301 19329 16313 19363
rect 16347 19360 16359 19363
rect 16574 19360 16580 19372
rect 16347 19332 16580 19360
rect 16347 19329 16359 19332
rect 16301 19323 16359 19329
rect 16316 19292 16344 19323
rect 16574 19320 16580 19332
rect 16632 19320 16638 19372
rect 16868 19369 16896 19400
rect 17512 19369 17540 19400
rect 19334 19388 19340 19400
rect 19392 19388 19398 19440
rect 19610 19388 19616 19440
rect 19668 19388 19674 19440
rect 22066 19375 22094 19468
rect 22296 19428 22324 19468
rect 22557 19465 22569 19499
rect 22603 19496 22615 19499
rect 22646 19496 22652 19508
rect 22603 19468 22652 19496
rect 22603 19465 22615 19468
rect 22557 19459 22615 19465
rect 22646 19456 22652 19468
rect 22704 19456 22710 19508
rect 22833 19431 22891 19437
rect 22833 19428 22845 19431
rect 22296 19400 22845 19428
rect 22833 19397 22845 19400
rect 22879 19397 22891 19431
rect 24210 19428 24216 19440
rect 24171 19400 24216 19428
rect 22833 19391 22891 19397
rect 24210 19388 24216 19400
rect 24268 19388 24274 19440
rect 17770 19369 17776 19372
rect 16853 19363 16911 19369
rect 16853 19329 16865 19363
rect 16899 19329 16911 19363
rect 16853 19323 16911 19329
rect 17129 19363 17187 19369
rect 17129 19329 17141 19363
rect 17175 19329 17187 19363
rect 17129 19323 17187 19329
rect 17497 19363 17555 19369
rect 17497 19329 17509 19363
rect 17543 19329 17555 19363
rect 17497 19323 17555 19329
rect 17764 19323 17776 19369
rect 17828 19360 17834 19372
rect 17828 19332 17864 19360
rect 15580 19264 16344 19292
rect 16592 19292 16620 19320
rect 17144 19292 17172 19323
rect 17770 19320 17776 19323
rect 17828 19320 17834 19332
rect 20070 19320 20076 19372
rect 20128 19360 20134 19372
rect 20358 19363 20416 19369
rect 20358 19360 20370 19363
rect 20128 19332 20370 19360
rect 20128 19320 20134 19332
rect 20358 19329 20370 19332
rect 20404 19329 20416 19363
rect 20622 19360 20628 19372
rect 20583 19332 20628 19360
rect 20358 19323 20416 19329
rect 20622 19320 20628 19332
rect 20680 19320 20686 19372
rect 20806 19320 20812 19372
rect 20864 19360 20870 19372
rect 21085 19363 21143 19369
rect 21085 19360 21097 19363
rect 20864 19332 21097 19360
rect 20864 19320 20870 19332
rect 21085 19329 21097 19332
rect 21131 19329 21143 19363
rect 21085 19323 21143 19329
rect 21269 19363 21327 19369
rect 21269 19329 21281 19363
rect 21315 19360 21327 19363
rect 21726 19360 21732 19372
rect 21315 19332 21732 19360
rect 21315 19329 21327 19332
rect 21269 19323 21327 19329
rect 21726 19320 21732 19332
rect 21784 19320 21790 19372
rect 22066 19369 22134 19375
rect 21913 19363 21971 19369
rect 21913 19329 21925 19363
rect 21959 19329 21971 19363
rect 22066 19338 22088 19369
rect 22076 19335 22088 19338
rect 22122 19335 22134 19369
rect 22076 19329 22134 19335
rect 22189 19363 22247 19369
rect 22189 19329 22201 19363
rect 22235 19329 22247 19363
rect 21913 19323 21971 19329
rect 22189 19323 22247 19329
rect 16592 19264 17172 19292
rect 14737 19255 14795 19261
rect 20898 19252 20904 19304
rect 20956 19292 20962 19304
rect 21928 19292 21956 19323
rect 20956 19264 21956 19292
rect 22204 19292 22232 19323
rect 22298 19320 22304 19372
rect 22356 19360 22362 19372
rect 23014 19360 23020 19372
rect 22356 19332 22401 19360
rect 22975 19332 23020 19360
rect 22356 19320 22362 19332
rect 23014 19320 23020 19332
rect 23072 19320 23078 19372
rect 23201 19363 23259 19369
rect 23201 19329 23213 19363
rect 23247 19360 23259 19363
rect 23290 19360 23296 19372
rect 23247 19332 23296 19360
rect 23247 19329 23259 19332
rect 23201 19323 23259 19329
rect 23290 19320 23296 19332
rect 23348 19360 23354 19372
rect 23477 19363 23535 19369
rect 23477 19360 23489 19363
rect 23348 19332 23489 19360
rect 23348 19320 23354 19332
rect 23477 19329 23489 19332
rect 23523 19329 23535 19363
rect 23658 19360 23664 19372
rect 23619 19332 23664 19360
rect 23477 19323 23535 19329
rect 23658 19320 23664 19332
rect 23716 19320 23722 19372
rect 22646 19292 22652 19304
rect 22204 19264 22652 19292
rect 20956 19252 20962 19264
rect 22646 19252 22652 19264
rect 22704 19252 22710 19304
rect 23566 19252 23572 19304
rect 23624 19292 23630 19304
rect 24670 19292 24676 19304
rect 23624 19264 24676 19292
rect 23624 19252 23630 19264
rect 24670 19252 24676 19264
rect 24728 19252 24734 19304
rect 11330 19224 11336 19236
rect 6886 19196 9904 19224
rect 9968 19196 11336 19224
rect 1578 19116 1584 19168
rect 1636 19156 1642 19168
rect 6886 19156 6914 19196
rect 1636 19128 6914 19156
rect 9876 19156 9904 19196
rect 11330 19184 11336 19196
rect 11388 19184 11394 19236
rect 14090 19184 14096 19236
rect 14148 19224 14154 19236
rect 15841 19227 15899 19233
rect 15841 19224 15853 19227
rect 14148 19196 15853 19224
rect 14148 19184 14154 19196
rect 15841 19193 15853 19196
rect 15887 19193 15899 19227
rect 15841 19187 15899 19193
rect 18432 19196 19748 19224
rect 14734 19156 14740 19168
rect 9876 19128 14740 19156
rect 1636 19116 1642 19128
rect 14734 19116 14740 19128
rect 14792 19116 14798 19168
rect 15105 19159 15163 19165
rect 15105 19125 15117 19159
rect 15151 19156 15163 19159
rect 15286 19156 15292 19168
rect 15151 19128 15292 19156
rect 15151 19125 15163 19128
rect 15105 19119 15163 19125
rect 15286 19116 15292 19128
rect 15344 19116 15350 19168
rect 15930 19116 15936 19168
rect 15988 19156 15994 19168
rect 16669 19159 16727 19165
rect 16669 19156 16681 19159
rect 15988 19128 16681 19156
rect 15988 19116 15994 19128
rect 16669 19125 16681 19128
rect 16715 19125 16727 19159
rect 16669 19119 16727 19125
rect 16758 19116 16764 19168
rect 16816 19156 16822 19168
rect 18432 19156 18460 19196
rect 16816 19128 18460 19156
rect 19245 19159 19303 19165
rect 16816 19116 16822 19128
rect 19245 19125 19257 19159
rect 19291 19156 19303 19159
rect 19610 19156 19616 19168
rect 19291 19128 19616 19156
rect 19291 19125 19303 19128
rect 19245 19119 19303 19125
rect 19610 19116 19616 19128
rect 19668 19116 19674 19168
rect 19720 19156 19748 19196
rect 23198 19184 23204 19236
rect 23256 19224 23262 19236
rect 23256 19196 23980 19224
rect 23256 19184 23262 19196
rect 23952 19168 23980 19196
rect 20714 19156 20720 19168
rect 19720 19128 20720 19156
rect 20714 19116 20720 19128
rect 20772 19116 20778 19168
rect 21450 19156 21456 19168
rect 21411 19128 21456 19156
rect 21450 19116 21456 19128
rect 21508 19116 21514 19168
rect 23842 19156 23848 19168
rect 23803 19128 23848 19156
rect 23842 19116 23848 19128
rect 23900 19116 23906 19168
rect 23934 19116 23940 19168
rect 23992 19156 23998 19168
rect 24305 19159 24363 19165
rect 24305 19156 24317 19159
rect 23992 19128 24317 19156
rect 23992 19116 23998 19128
rect 24305 19125 24317 19128
rect 24351 19125 24363 19159
rect 24305 19119 24363 19125
rect 1104 19066 28888 19088
rect 1104 19014 5582 19066
rect 5634 19014 5646 19066
rect 5698 19014 5710 19066
rect 5762 19014 5774 19066
rect 5826 19014 5838 19066
rect 5890 19014 14846 19066
rect 14898 19014 14910 19066
rect 14962 19014 14974 19066
rect 15026 19014 15038 19066
rect 15090 19014 15102 19066
rect 15154 19014 24110 19066
rect 24162 19014 24174 19066
rect 24226 19014 24238 19066
rect 24290 19014 24302 19066
rect 24354 19014 24366 19066
rect 24418 19014 28888 19066
rect 1104 18992 28888 19014
rect 8846 18912 8852 18964
rect 8904 18952 8910 18964
rect 8941 18955 8999 18961
rect 8941 18952 8953 18955
rect 8904 18924 8953 18952
rect 8904 18912 8910 18924
rect 8941 18921 8953 18924
rect 8987 18921 8999 18955
rect 8941 18915 8999 18921
rect 10870 18912 10876 18964
rect 10928 18952 10934 18964
rect 12437 18955 12495 18961
rect 10928 18924 11192 18952
rect 10928 18912 10934 18924
rect 7668 18856 11100 18884
rect 1394 18748 1400 18760
rect 1355 18720 1400 18748
rect 1394 18708 1400 18720
rect 1452 18708 1458 18760
rect 6638 18748 6644 18760
rect 6599 18720 6644 18748
rect 6638 18708 6644 18720
rect 6696 18708 6702 18760
rect 6914 18757 6920 18760
rect 6908 18711 6920 18757
rect 6972 18748 6978 18760
rect 6972 18720 7008 18748
rect 6914 18708 6920 18711
rect 6972 18708 6978 18720
rect 7282 18708 7288 18760
rect 7340 18748 7346 18760
rect 7668 18748 7696 18856
rect 8110 18776 8116 18828
rect 8168 18816 8174 18828
rect 9493 18819 9551 18825
rect 9493 18816 9505 18819
rect 8168 18788 9505 18816
rect 8168 18776 8174 18788
rect 9493 18785 9505 18788
rect 9539 18785 9551 18819
rect 10962 18816 10968 18828
rect 10923 18788 10968 18816
rect 9493 18779 9551 18785
rect 10962 18776 10968 18788
rect 11020 18776 11026 18828
rect 7340 18720 7696 18748
rect 9309 18751 9367 18757
rect 7340 18708 7346 18720
rect 9309 18717 9321 18751
rect 9355 18748 9367 18751
rect 9674 18748 9680 18760
rect 9355 18720 9680 18748
rect 9355 18717 9367 18720
rect 9309 18711 9367 18717
rect 9674 18708 9680 18720
rect 9732 18748 9738 18760
rect 10873 18751 10931 18757
rect 10873 18748 10885 18751
rect 9732 18720 10885 18748
rect 9732 18708 9738 18720
rect 10873 18717 10885 18720
rect 10919 18717 10931 18751
rect 10873 18711 10931 18717
rect 9401 18683 9459 18689
rect 9401 18680 9413 18683
rect 8036 18652 9413 18680
rect 7834 18572 7840 18624
rect 7892 18612 7898 18624
rect 8036 18621 8064 18652
rect 9401 18649 9413 18652
rect 9447 18680 9459 18683
rect 9582 18680 9588 18692
rect 9447 18652 9588 18680
rect 9447 18649 9459 18652
rect 9401 18643 9459 18649
rect 9582 18640 9588 18652
rect 9640 18640 9646 18692
rect 11072 18680 11100 18856
rect 11164 18748 11192 18924
rect 12437 18921 12449 18955
rect 12483 18952 12495 18955
rect 12710 18952 12716 18964
rect 12483 18924 12716 18952
rect 12483 18921 12495 18924
rect 12437 18915 12495 18921
rect 12710 18912 12716 18924
rect 12768 18952 12774 18964
rect 13081 18955 13139 18961
rect 13081 18952 13093 18955
rect 12768 18924 13093 18952
rect 12768 18912 12774 18924
rect 13081 18921 13093 18924
rect 13127 18921 13139 18955
rect 13081 18915 13139 18921
rect 14366 18912 14372 18964
rect 14424 18952 14430 18964
rect 16758 18952 16764 18964
rect 14424 18924 16764 18952
rect 14424 18912 14430 18924
rect 16758 18912 16764 18924
rect 16816 18912 16822 18964
rect 17770 18912 17776 18964
rect 17828 18952 17834 18964
rect 17865 18955 17923 18961
rect 17865 18952 17877 18955
rect 17828 18924 17877 18952
rect 17828 18912 17834 18924
rect 17865 18921 17877 18924
rect 17911 18921 17923 18955
rect 17865 18915 17923 18921
rect 18693 18955 18751 18961
rect 18693 18921 18705 18955
rect 18739 18952 18751 18955
rect 19334 18952 19340 18964
rect 18739 18924 19340 18952
rect 18739 18921 18751 18924
rect 18693 18915 18751 18921
rect 19334 18912 19340 18924
rect 19392 18952 19398 18964
rect 20622 18952 20628 18964
rect 19392 18924 20628 18952
rect 19392 18912 19398 18924
rect 20622 18912 20628 18924
rect 20680 18912 20686 18964
rect 20714 18912 20720 18964
rect 20772 18952 20778 18964
rect 21913 18955 21971 18961
rect 20772 18924 21680 18952
rect 20772 18912 20778 18924
rect 13814 18844 13820 18896
rect 13872 18884 13878 18896
rect 13872 18856 14504 18884
rect 13872 18844 13878 18856
rect 14093 18819 14151 18825
rect 14093 18816 14105 18819
rect 11532 18788 14105 18816
rect 11425 18751 11483 18757
rect 11425 18748 11437 18751
rect 11164 18720 11437 18748
rect 11425 18717 11437 18720
rect 11471 18717 11483 18751
rect 11425 18711 11483 18717
rect 11532 18680 11560 18788
rect 14093 18785 14105 18788
rect 14139 18785 14151 18819
rect 14093 18779 14151 18785
rect 12544 18720 13140 18748
rect 12250 18680 12256 18692
rect 11072 18652 11560 18680
rect 12211 18652 12256 18680
rect 12250 18640 12256 18652
rect 12308 18640 12314 18692
rect 8021 18615 8079 18621
rect 8021 18612 8033 18615
rect 7892 18584 8033 18612
rect 7892 18572 7898 18584
rect 8021 18581 8033 18584
rect 8067 18581 8079 18615
rect 8021 18575 8079 18581
rect 10413 18615 10471 18621
rect 10413 18581 10425 18615
rect 10459 18612 10471 18615
rect 10686 18612 10692 18624
rect 10459 18584 10692 18612
rect 10459 18581 10471 18584
rect 10413 18575 10471 18581
rect 10686 18572 10692 18584
rect 10744 18572 10750 18624
rect 10781 18615 10839 18621
rect 10781 18581 10793 18615
rect 10827 18612 10839 18615
rect 11422 18612 11428 18624
rect 10827 18584 11428 18612
rect 10827 18581 10839 18584
rect 10781 18575 10839 18581
rect 11422 18572 11428 18584
rect 11480 18572 11486 18624
rect 11606 18612 11612 18624
rect 11567 18584 11612 18612
rect 11606 18572 11612 18584
rect 11664 18572 11670 18624
rect 12434 18572 12440 18624
rect 12492 18621 12498 18624
rect 12492 18615 12511 18621
rect 12499 18612 12511 18615
rect 12544 18612 12572 18720
rect 12802 18640 12808 18692
rect 12860 18680 12866 18692
rect 13112 18689 13140 18720
rect 14182 18708 14188 18760
rect 14240 18748 14246 18760
rect 14366 18748 14372 18760
rect 14240 18720 14372 18748
rect 14240 18708 14246 18720
rect 14366 18708 14372 18720
rect 14424 18708 14430 18760
rect 14476 18757 14504 18856
rect 14550 18844 14556 18896
rect 14608 18844 14614 18896
rect 14734 18844 14740 18896
rect 14792 18884 14798 18896
rect 15565 18887 15623 18893
rect 14792 18856 15516 18884
rect 14792 18844 14798 18856
rect 14568 18816 14596 18844
rect 15102 18816 15108 18828
rect 14568 18788 14780 18816
rect 15063 18788 15108 18816
rect 14458 18751 14516 18757
rect 14458 18717 14470 18751
rect 14504 18717 14516 18751
rect 14458 18711 14516 18717
rect 14553 18751 14611 18757
rect 14553 18717 14565 18751
rect 14599 18748 14611 18751
rect 14642 18748 14648 18760
rect 14599 18720 14648 18748
rect 14599 18717 14611 18720
rect 14553 18711 14611 18717
rect 14642 18708 14648 18720
rect 14700 18708 14706 18760
rect 14752 18757 14780 18788
rect 15102 18776 15108 18788
rect 15160 18776 15166 18828
rect 15488 18816 15516 18856
rect 15565 18853 15577 18887
rect 15611 18884 15623 18887
rect 15611 18856 21588 18884
rect 15611 18853 15623 18856
rect 15565 18847 15623 18853
rect 17310 18816 17316 18828
rect 15488 18788 17316 18816
rect 17310 18776 17316 18788
rect 17368 18776 17374 18828
rect 17770 18816 17776 18828
rect 17512 18788 17776 18816
rect 14737 18751 14795 18757
rect 14737 18717 14749 18751
rect 14783 18717 14795 18751
rect 14737 18711 14795 18717
rect 14826 18708 14832 18760
rect 14884 18748 14890 18760
rect 15013 18751 15071 18757
rect 15013 18748 15025 18751
rect 14884 18720 15025 18748
rect 14884 18708 14890 18720
rect 15013 18717 15025 18720
rect 15059 18717 15071 18751
rect 15286 18748 15292 18760
rect 15247 18720 15292 18748
rect 15013 18711 15071 18717
rect 15286 18708 15292 18720
rect 15344 18708 15350 18760
rect 15381 18751 15439 18757
rect 15381 18717 15393 18751
rect 15427 18717 15439 18751
rect 15381 18711 15439 18717
rect 12897 18683 12955 18689
rect 12897 18680 12909 18683
rect 12860 18652 12909 18680
rect 12860 18640 12866 18652
rect 12897 18649 12909 18652
rect 12943 18649 12955 18683
rect 12897 18643 12955 18649
rect 13097 18683 13155 18689
rect 13097 18649 13109 18683
rect 13143 18649 13155 18683
rect 13097 18643 13155 18649
rect 13188 18652 14412 18680
rect 12499 18584 12572 18612
rect 12621 18615 12679 18621
rect 12499 18581 12511 18584
rect 12492 18575 12511 18581
rect 12621 18581 12633 18615
rect 12667 18612 12679 18615
rect 13188 18612 13216 18652
rect 12667 18584 13216 18612
rect 13265 18615 13323 18621
rect 12667 18581 12679 18584
rect 12621 18575 12679 18581
rect 13265 18581 13277 18615
rect 13311 18612 13323 18615
rect 13998 18612 14004 18624
rect 13311 18584 14004 18612
rect 13311 18581 13323 18584
rect 13265 18575 13323 18581
rect 12492 18572 12498 18575
rect 13998 18572 14004 18584
rect 14056 18572 14062 18624
rect 14384 18612 14412 18652
rect 15396 18612 15424 18711
rect 16022 18708 16028 18760
rect 16080 18748 16086 18760
rect 16117 18751 16175 18757
rect 16117 18748 16129 18751
rect 16080 18720 16129 18748
rect 16080 18708 16086 18720
rect 16117 18717 16129 18720
rect 16163 18717 16175 18751
rect 16117 18711 16175 18717
rect 16393 18751 16451 18757
rect 16393 18717 16405 18751
rect 16439 18748 16451 18751
rect 16574 18748 16580 18760
rect 16439 18720 16580 18748
rect 16439 18717 16451 18720
rect 16393 18711 16451 18717
rect 16574 18708 16580 18720
rect 16632 18748 16638 18760
rect 16942 18748 16948 18760
rect 16632 18720 16948 18748
rect 16632 18708 16638 18720
rect 16942 18708 16948 18720
rect 17000 18708 17006 18760
rect 17221 18751 17279 18757
rect 17221 18717 17233 18751
rect 17267 18717 17279 18751
rect 17402 18748 17408 18760
rect 17363 18720 17408 18748
rect 17221 18711 17279 18717
rect 16301 18683 16359 18689
rect 16301 18649 16313 18683
rect 16347 18680 16359 18683
rect 16666 18680 16672 18692
rect 16347 18652 16672 18680
rect 16347 18649 16359 18652
rect 16301 18643 16359 18649
rect 16666 18640 16672 18652
rect 16724 18640 16730 18692
rect 17236 18680 17264 18711
rect 17402 18708 17408 18720
rect 17460 18708 17466 18760
rect 17512 18757 17540 18788
rect 17770 18776 17776 18788
rect 17828 18776 17834 18828
rect 19429 18819 19487 18825
rect 19429 18785 19441 18819
rect 19475 18816 19487 18819
rect 19475 18788 20576 18816
rect 19475 18785 19487 18788
rect 19429 18779 19487 18785
rect 17497 18751 17555 18757
rect 17497 18717 17509 18751
rect 17543 18717 17555 18751
rect 17497 18711 17555 18717
rect 17589 18751 17647 18757
rect 17589 18717 17601 18751
rect 17635 18748 17647 18751
rect 17678 18748 17684 18760
rect 17635 18720 17684 18748
rect 17635 18717 17647 18720
rect 17589 18711 17647 18717
rect 17678 18708 17684 18720
rect 17736 18748 17742 18760
rect 17954 18748 17960 18760
rect 17736 18720 17960 18748
rect 17736 18708 17742 18720
rect 17954 18708 17960 18720
rect 18012 18708 18018 18760
rect 18138 18748 18144 18760
rect 18099 18720 18144 18748
rect 18138 18708 18144 18720
rect 18196 18708 18202 18760
rect 18785 18751 18843 18757
rect 18785 18717 18797 18751
rect 18831 18748 18843 18751
rect 20254 18748 20260 18760
rect 18831 18720 20260 18748
rect 18831 18717 18843 18720
rect 18785 18711 18843 18717
rect 20254 18708 20260 18720
rect 20312 18708 20318 18760
rect 20548 18757 20576 18788
rect 20349 18751 20407 18757
rect 20349 18717 20361 18751
rect 20395 18717 20407 18751
rect 20349 18711 20407 18717
rect 20441 18751 20499 18757
rect 20441 18717 20453 18751
rect 20487 18717 20499 18751
rect 20441 18711 20499 18717
rect 20533 18751 20591 18757
rect 20533 18717 20545 18751
rect 20579 18717 20591 18751
rect 20714 18748 20720 18760
rect 20675 18720 20720 18748
rect 20533 18711 20591 18717
rect 19242 18680 19248 18692
rect 16868 18652 19248 18680
rect 14384 18584 15424 18612
rect 15654 18572 15660 18624
rect 15712 18612 15718 18624
rect 15933 18615 15991 18621
rect 15933 18612 15945 18615
rect 15712 18584 15945 18612
rect 15712 18572 15718 18584
rect 15933 18581 15945 18584
rect 15979 18581 15991 18615
rect 15933 18575 15991 18581
rect 16206 18572 16212 18624
rect 16264 18612 16270 18624
rect 16868 18612 16896 18652
rect 19242 18640 19248 18652
rect 19300 18640 19306 18692
rect 19610 18680 19616 18692
rect 19571 18652 19616 18680
rect 19610 18640 19616 18652
rect 19668 18640 19674 18692
rect 19797 18683 19855 18689
rect 19797 18649 19809 18683
rect 19843 18680 19855 18683
rect 20162 18680 20168 18692
rect 19843 18652 20168 18680
rect 19843 18649 19855 18652
rect 19797 18643 19855 18649
rect 20162 18640 20168 18652
rect 20220 18640 20226 18692
rect 16264 18584 16896 18612
rect 16945 18615 17003 18621
rect 16264 18572 16270 18584
rect 16945 18581 16957 18615
rect 16991 18612 17003 18615
rect 18046 18612 18052 18624
rect 16991 18584 18052 18612
rect 16991 18581 17003 18584
rect 16945 18575 17003 18581
rect 18046 18572 18052 18584
rect 18104 18572 18110 18624
rect 18322 18612 18328 18624
rect 18283 18584 18328 18612
rect 18322 18572 18328 18584
rect 18380 18572 18386 18624
rect 20070 18612 20076 18624
rect 20031 18584 20076 18612
rect 20070 18572 20076 18584
rect 20128 18572 20134 18624
rect 20364 18612 20392 18711
rect 20456 18680 20484 18711
rect 20714 18708 20720 18720
rect 20772 18708 20778 18760
rect 21174 18708 21180 18760
rect 21232 18748 21238 18760
rect 21269 18751 21327 18757
rect 21269 18748 21281 18751
rect 21232 18720 21281 18748
rect 21232 18708 21238 18720
rect 21269 18717 21281 18720
rect 21315 18717 21327 18751
rect 21450 18748 21456 18760
rect 21411 18720 21456 18748
rect 21269 18711 21327 18717
rect 20622 18680 20628 18692
rect 20456 18652 20628 18680
rect 20622 18640 20628 18652
rect 20680 18640 20686 18692
rect 20530 18612 20536 18624
rect 20364 18584 20536 18612
rect 20530 18572 20536 18584
rect 20588 18572 20594 18624
rect 21284 18612 21312 18711
rect 21450 18708 21456 18720
rect 21508 18708 21514 18760
rect 21560 18757 21588 18856
rect 21652 18757 21680 18924
rect 21913 18921 21925 18955
rect 21959 18952 21971 18955
rect 22370 18952 22376 18964
rect 21959 18924 22376 18952
rect 21959 18921 21971 18924
rect 21913 18915 21971 18921
rect 22370 18912 22376 18924
rect 22428 18912 22434 18964
rect 23658 18912 23664 18964
rect 23716 18952 23722 18964
rect 25777 18955 25835 18961
rect 25777 18952 25789 18955
rect 23716 18924 25789 18952
rect 23716 18912 23722 18924
rect 25777 18921 25789 18924
rect 25823 18921 25835 18955
rect 25777 18915 25835 18921
rect 21818 18844 21824 18896
rect 21876 18884 21882 18896
rect 22833 18887 22891 18893
rect 22833 18884 22845 18887
rect 21876 18856 22845 18884
rect 21876 18844 21882 18856
rect 22833 18853 22845 18856
rect 22879 18853 22891 18887
rect 23676 18884 23704 18912
rect 22833 18847 22891 18853
rect 22931 18856 23704 18884
rect 22931 18816 22959 18856
rect 23842 18816 23848 18828
rect 22388 18788 22959 18816
rect 23400 18788 23848 18816
rect 21545 18751 21603 18757
rect 21545 18717 21557 18751
rect 21591 18717 21603 18751
rect 21545 18711 21603 18717
rect 21637 18751 21695 18757
rect 21637 18717 21649 18751
rect 21683 18748 21695 18751
rect 22278 18748 22284 18760
rect 21683 18720 22284 18748
rect 21683 18717 21695 18720
rect 21637 18711 21695 18717
rect 22278 18708 22284 18720
rect 22336 18708 22342 18760
rect 22388 18757 22416 18788
rect 22373 18751 22431 18757
rect 22373 18717 22385 18751
rect 22419 18717 22431 18751
rect 22373 18711 22431 18717
rect 22922 18708 22928 18760
rect 22980 18748 22986 18760
rect 23400 18757 23428 18788
rect 23842 18776 23848 18788
rect 23900 18776 23906 18828
rect 23474 18757 23480 18760
rect 23201 18751 23259 18757
rect 23201 18748 23213 18751
rect 22980 18720 23213 18748
rect 22980 18708 22986 18720
rect 23201 18717 23213 18720
rect 23247 18717 23259 18751
rect 23201 18711 23259 18717
rect 23364 18751 23428 18757
rect 23364 18717 23376 18751
rect 23410 18720 23428 18751
rect 23464 18751 23480 18757
rect 23410 18717 23422 18720
rect 23364 18711 23422 18717
rect 23464 18717 23476 18751
rect 23464 18711 23480 18717
rect 23474 18708 23480 18711
rect 23532 18708 23538 18760
rect 23566 18708 23572 18760
rect 23624 18757 23630 18760
rect 23624 18751 23647 18757
rect 23635 18717 23647 18751
rect 23624 18711 23647 18717
rect 23624 18708 23630 18711
rect 23934 18708 23940 18760
rect 23992 18748 23998 18760
rect 24397 18751 24455 18757
rect 24397 18748 24409 18751
rect 23992 18720 24409 18748
rect 23992 18708 23998 18720
rect 24397 18717 24409 18720
rect 24443 18717 24455 18751
rect 24397 18711 24455 18717
rect 21726 18640 21732 18692
rect 21784 18680 21790 18692
rect 22189 18683 22247 18689
rect 22189 18680 22201 18683
rect 21784 18652 22201 18680
rect 21784 18640 21790 18652
rect 22189 18649 22201 18652
rect 22235 18649 22247 18683
rect 22189 18643 22247 18649
rect 23845 18683 23903 18689
rect 23845 18649 23857 18683
rect 23891 18680 23903 18683
rect 24642 18683 24700 18689
rect 24642 18680 24654 18683
rect 23891 18652 24654 18680
rect 23891 18649 23903 18652
rect 23845 18643 23903 18649
rect 24642 18649 24654 18652
rect 24688 18649 24700 18683
rect 24642 18643 24700 18649
rect 21818 18612 21824 18624
rect 21284 18584 21824 18612
rect 21818 18572 21824 18584
rect 21876 18572 21882 18624
rect 22002 18572 22008 18624
rect 22060 18612 22066 18624
rect 22557 18615 22615 18621
rect 22557 18612 22569 18615
rect 22060 18584 22569 18612
rect 22060 18572 22066 18584
rect 22557 18581 22569 18584
rect 22603 18581 22615 18615
rect 22557 18575 22615 18581
rect 22646 18572 22652 18624
rect 22704 18612 22710 18624
rect 23474 18612 23480 18624
rect 22704 18584 23480 18612
rect 22704 18572 22710 18584
rect 23474 18572 23480 18584
rect 23532 18572 23538 18624
rect 1104 18522 28888 18544
rect 1104 18470 10214 18522
rect 10266 18470 10278 18522
rect 10330 18470 10342 18522
rect 10394 18470 10406 18522
rect 10458 18470 10470 18522
rect 10522 18470 19478 18522
rect 19530 18470 19542 18522
rect 19594 18470 19606 18522
rect 19658 18470 19670 18522
rect 19722 18470 19734 18522
rect 19786 18470 28888 18522
rect 1104 18448 28888 18470
rect 7006 18368 7012 18420
rect 7064 18408 7070 18420
rect 7101 18411 7159 18417
rect 7101 18408 7113 18411
rect 7064 18380 7113 18408
rect 7064 18368 7070 18380
rect 7101 18377 7113 18380
rect 7147 18377 7159 18411
rect 7101 18371 7159 18377
rect 7469 18411 7527 18417
rect 7469 18377 7481 18411
rect 7515 18377 7527 18411
rect 7834 18408 7840 18420
rect 7795 18380 7840 18408
rect 7469 18371 7527 18377
rect 5741 18275 5799 18281
rect 5741 18241 5753 18275
rect 5787 18272 5799 18275
rect 6917 18275 6975 18281
rect 5787 18244 6868 18272
rect 5787 18241 5799 18244
rect 5741 18235 5799 18241
rect 5994 18204 6000 18216
rect 5955 18176 6000 18204
rect 5994 18164 6000 18176
rect 6052 18164 6058 18216
rect 6730 18204 6736 18216
rect 6691 18176 6736 18204
rect 6730 18164 6736 18176
rect 6788 18164 6794 18216
rect 6840 18204 6868 18244
rect 6917 18241 6929 18275
rect 6963 18272 6975 18275
rect 7484 18272 7512 18371
rect 7834 18368 7840 18380
rect 7892 18368 7898 18420
rect 8573 18411 8631 18417
rect 8573 18377 8585 18411
rect 8619 18408 8631 18411
rect 9030 18408 9036 18420
rect 8619 18380 9036 18408
rect 8619 18377 8631 18380
rect 8573 18371 8631 18377
rect 6963 18244 7512 18272
rect 6963 18241 6975 18244
rect 6917 18235 6975 18241
rect 7282 18204 7288 18216
rect 6840 18176 7288 18204
rect 7282 18164 7288 18176
rect 7340 18164 7346 18216
rect 7374 18164 7380 18216
rect 7432 18204 7438 18216
rect 7929 18207 7987 18213
rect 7929 18204 7941 18207
rect 7432 18176 7941 18204
rect 7432 18164 7438 18176
rect 7929 18173 7941 18176
rect 7975 18173 7987 18207
rect 8110 18204 8116 18216
rect 8071 18176 8116 18204
rect 7929 18167 7987 18173
rect 8110 18164 8116 18176
rect 8168 18164 8174 18216
rect 6012 18136 6040 18164
rect 6638 18136 6644 18148
rect 6012 18108 6644 18136
rect 6638 18096 6644 18108
rect 6696 18136 6702 18148
rect 8588 18136 8616 18371
rect 9030 18368 9036 18380
rect 9088 18368 9094 18420
rect 9582 18408 9588 18420
rect 9543 18380 9588 18408
rect 9582 18368 9588 18380
rect 9640 18368 9646 18420
rect 9674 18368 9680 18420
rect 9732 18408 9738 18420
rect 10962 18408 10968 18420
rect 9732 18380 10968 18408
rect 9732 18368 9738 18380
rect 10962 18368 10968 18380
rect 11020 18368 11026 18420
rect 11422 18368 11428 18420
rect 11480 18408 11486 18420
rect 12897 18411 12955 18417
rect 12897 18408 12909 18411
rect 11480 18380 12909 18408
rect 11480 18368 11486 18380
rect 12897 18377 12909 18380
rect 12943 18408 12955 18411
rect 13814 18408 13820 18420
rect 12943 18380 13216 18408
rect 13775 18380 13820 18408
rect 12943 18377 12955 18380
rect 12897 18371 12955 18377
rect 8665 18343 8723 18349
rect 8665 18309 8677 18343
rect 8711 18340 8723 18343
rect 9858 18340 9864 18352
rect 8711 18312 9864 18340
rect 8711 18309 8723 18312
rect 8665 18303 8723 18309
rect 9858 18300 9864 18312
rect 9916 18300 9922 18352
rect 13078 18340 13084 18352
rect 10520 18312 13084 18340
rect 9493 18275 9551 18281
rect 9493 18241 9505 18275
rect 9539 18272 9551 18275
rect 10318 18272 10324 18284
rect 9539 18244 10324 18272
rect 9539 18241 9551 18244
rect 9493 18235 9551 18241
rect 10318 18232 10324 18244
rect 10376 18232 10382 18284
rect 9674 18204 9680 18216
rect 9635 18176 9680 18204
rect 9674 18164 9680 18176
rect 9732 18164 9738 18216
rect 9766 18164 9772 18216
rect 9824 18204 9830 18216
rect 10413 18207 10471 18213
rect 10413 18204 10425 18207
rect 9824 18176 10425 18204
rect 9824 18164 9830 18176
rect 10413 18173 10425 18176
rect 10459 18173 10471 18207
rect 10413 18167 10471 18173
rect 6696 18108 8616 18136
rect 8956 18108 9628 18136
rect 6696 18096 6702 18108
rect 4614 18068 4620 18080
rect 4575 18040 4620 18068
rect 4614 18028 4620 18040
rect 4672 18028 4678 18080
rect 6730 18028 6736 18080
rect 6788 18068 6794 18080
rect 8956 18068 8984 18108
rect 9122 18068 9128 18080
rect 6788 18040 8984 18068
rect 9083 18040 9128 18068
rect 6788 18028 6794 18040
rect 9122 18028 9128 18040
rect 9180 18028 9186 18080
rect 9600 18068 9628 18108
rect 10520 18068 10548 18312
rect 13078 18300 13084 18312
rect 13136 18300 13142 18352
rect 13188 18349 13216 18380
rect 13814 18368 13820 18380
rect 13872 18368 13878 18420
rect 14642 18368 14648 18420
rect 14700 18408 14706 18420
rect 19613 18411 19671 18417
rect 14700 18380 19472 18408
rect 14700 18368 14706 18380
rect 13173 18343 13231 18349
rect 13173 18309 13185 18343
rect 13219 18309 13231 18343
rect 13173 18303 13231 18309
rect 13389 18343 13447 18349
rect 13389 18309 13401 18343
rect 13435 18340 13447 18343
rect 13538 18340 13544 18352
rect 13435 18312 13544 18340
rect 13435 18309 13447 18312
rect 13389 18303 13447 18309
rect 13538 18300 13544 18312
rect 13596 18300 13602 18352
rect 15746 18340 15752 18352
rect 14936 18312 15752 18340
rect 10597 18275 10655 18281
rect 10597 18241 10609 18275
rect 10643 18272 10655 18275
rect 10686 18272 10692 18284
rect 10643 18244 10692 18272
rect 10643 18241 10655 18244
rect 10597 18235 10655 18241
rect 10686 18232 10692 18244
rect 10744 18232 10750 18284
rect 11146 18232 11152 18284
rect 11204 18272 11210 18284
rect 11773 18275 11831 18281
rect 11773 18272 11785 18275
rect 11204 18244 11785 18272
rect 11204 18232 11210 18244
rect 11773 18241 11785 18244
rect 11819 18241 11831 18275
rect 13998 18272 14004 18284
rect 13959 18244 14004 18272
rect 11773 18235 11831 18241
rect 13998 18232 14004 18244
rect 14056 18232 14062 18284
rect 14090 18232 14096 18284
rect 14148 18272 14154 18284
rect 14366 18272 14372 18284
rect 14148 18244 14193 18272
rect 14327 18244 14372 18272
rect 14148 18232 14154 18244
rect 14366 18232 14372 18244
rect 14424 18232 14430 18284
rect 14936 18281 14964 18312
rect 15746 18300 15752 18312
rect 15804 18300 15810 18352
rect 17034 18300 17040 18352
rect 17092 18340 17098 18352
rect 17310 18340 17316 18352
rect 17092 18312 17316 18340
rect 17092 18300 17098 18312
rect 17310 18300 17316 18312
rect 17368 18340 17374 18352
rect 17773 18343 17831 18349
rect 17773 18340 17785 18343
rect 17368 18312 17785 18340
rect 17368 18300 17374 18312
rect 17773 18309 17785 18312
rect 17819 18309 17831 18343
rect 19334 18340 19340 18352
rect 17773 18303 17831 18309
rect 18248 18312 19340 18340
rect 14829 18275 14887 18281
rect 14829 18241 14841 18275
rect 14875 18241 14887 18275
rect 14829 18235 14887 18241
rect 14921 18275 14979 18281
rect 14921 18241 14933 18275
rect 14967 18241 14979 18275
rect 14921 18235 14979 18241
rect 15197 18275 15255 18281
rect 15197 18241 15209 18275
rect 15243 18272 15255 18275
rect 15286 18272 15292 18284
rect 15243 18244 15292 18272
rect 15243 18241 15255 18244
rect 15197 18235 15255 18241
rect 11514 18204 11520 18216
rect 11475 18176 11520 18204
rect 11514 18164 11520 18176
rect 11572 18164 11578 18216
rect 14844 18204 14872 18235
rect 15286 18232 15292 18244
rect 15344 18232 15350 18284
rect 16022 18272 16028 18284
rect 15983 18244 16028 18272
rect 16022 18232 16028 18244
rect 16080 18232 16086 18284
rect 16942 18272 16948 18284
rect 16903 18244 16948 18272
rect 16942 18232 16948 18244
rect 17000 18232 17006 18284
rect 18248 18281 18276 18312
rect 19334 18300 19340 18312
rect 19392 18300 19398 18352
rect 19444 18340 19472 18380
rect 19613 18377 19625 18411
rect 19659 18408 19671 18411
rect 19886 18408 19892 18420
rect 19659 18380 19892 18408
rect 19659 18377 19671 18380
rect 19613 18371 19671 18377
rect 19886 18368 19892 18380
rect 19944 18368 19950 18420
rect 20162 18368 20168 18420
rect 20220 18408 20226 18420
rect 20220 18380 21312 18408
rect 20220 18368 20226 18380
rect 20257 18343 20315 18349
rect 20257 18340 20269 18343
rect 19444 18312 20269 18340
rect 20257 18309 20269 18312
rect 20303 18309 20315 18343
rect 20438 18340 20444 18352
rect 20399 18312 20444 18340
rect 20257 18303 20315 18309
rect 20438 18300 20444 18312
rect 20496 18300 20502 18352
rect 20714 18340 20720 18352
rect 20548 18312 20720 18340
rect 18233 18275 18291 18281
rect 18233 18241 18245 18275
rect 18279 18241 18291 18275
rect 18233 18235 18291 18241
rect 18322 18232 18328 18284
rect 18380 18272 18386 18284
rect 18489 18275 18547 18281
rect 18489 18272 18501 18275
rect 18380 18244 18501 18272
rect 18380 18232 18386 18244
rect 18489 18241 18501 18244
rect 18535 18241 18547 18275
rect 18489 18235 18547 18241
rect 19242 18232 19248 18284
rect 19300 18272 19306 18284
rect 20548 18272 20576 18312
rect 20714 18300 20720 18312
rect 20772 18340 20778 18352
rect 20898 18340 20904 18352
rect 20772 18312 20904 18340
rect 20772 18300 20778 18312
rect 20898 18300 20904 18312
rect 20956 18300 20962 18352
rect 21284 18349 21312 18380
rect 22094 18368 22100 18420
rect 22152 18368 22158 18420
rect 22462 18408 22468 18420
rect 22423 18380 22468 18408
rect 22462 18368 22468 18380
rect 22520 18368 22526 18420
rect 21269 18343 21327 18349
rect 21269 18309 21281 18343
rect 21315 18340 21327 18343
rect 21910 18340 21916 18352
rect 21315 18312 21916 18340
rect 21315 18309 21327 18312
rect 21269 18303 21327 18309
rect 21910 18300 21916 18312
rect 21968 18300 21974 18352
rect 19300 18244 20576 18272
rect 20625 18275 20683 18281
rect 19300 18232 19306 18244
rect 20625 18241 20637 18275
rect 20671 18272 20683 18275
rect 20806 18272 20812 18284
rect 20671 18244 20812 18272
rect 20671 18241 20683 18244
rect 20625 18235 20683 18241
rect 20806 18232 20812 18244
rect 20864 18232 20870 18284
rect 21082 18272 21088 18284
rect 21043 18244 21088 18272
rect 21082 18232 21088 18244
rect 21140 18232 21146 18284
rect 21818 18272 21824 18284
rect 21779 18244 21824 18272
rect 21818 18232 21824 18244
rect 21876 18232 21882 18284
rect 22002 18272 22008 18284
rect 21963 18244 22008 18272
rect 22002 18232 22008 18244
rect 22060 18232 22066 18284
rect 22112 18281 22140 18368
rect 22738 18300 22744 18352
rect 22796 18340 22802 18352
rect 23477 18343 23535 18349
rect 22796 18312 23264 18340
rect 22796 18300 22802 18312
rect 22097 18275 22155 18281
rect 22097 18241 22109 18275
rect 22143 18241 22155 18275
rect 22097 18235 22155 18241
rect 22189 18275 22247 18281
rect 22189 18241 22201 18275
rect 22235 18272 22247 18275
rect 22278 18272 22284 18284
rect 22235 18244 22284 18272
rect 22235 18241 22247 18244
rect 22189 18235 22247 18241
rect 22278 18232 22284 18244
rect 22336 18232 22342 18284
rect 23014 18281 23020 18284
rect 22833 18275 22891 18281
rect 22833 18241 22845 18275
rect 22879 18241 22891 18275
rect 23012 18272 23020 18281
rect 22975 18244 23020 18272
rect 22833 18235 22891 18241
rect 23012 18235 23020 18244
rect 15102 18204 15108 18216
rect 13556 18176 14872 18204
rect 15015 18176 15108 18204
rect 13556 18145 13584 18176
rect 13541 18139 13599 18145
rect 13541 18105 13553 18139
rect 13587 18105 13599 18139
rect 13541 18099 13599 18105
rect 14277 18139 14335 18145
rect 14277 18105 14289 18139
rect 14323 18136 14335 18139
rect 15028 18136 15056 18176
rect 15102 18164 15108 18176
rect 15160 18204 15166 18216
rect 15470 18204 15476 18216
rect 15160 18176 15476 18204
rect 15160 18164 15166 18176
rect 15470 18164 15476 18176
rect 15528 18164 15534 18216
rect 16301 18207 16359 18213
rect 16301 18173 16313 18207
rect 16347 18204 16359 18207
rect 16390 18204 16396 18216
rect 16347 18176 16396 18204
rect 16347 18173 16359 18176
rect 16301 18167 16359 18173
rect 16390 18164 16396 18176
rect 16448 18164 16454 18216
rect 16666 18204 16672 18216
rect 16627 18176 16672 18204
rect 16666 18164 16672 18176
rect 16724 18164 16730 18216
rect 20530 18136 20536 18148
rect 14323 18108 15056 18136
rect 19904 18108 20536 18136
rect 14323 18105 14335 18108
rect 14277 18099 14335 18105
rect 9600 18040 10548 18068
rect 10781 18071 10839 18077
rect 10781 18037 10793 18071
rect 10827 18068 10839 18071
rect 10962 18068 10968 18080
rect 10827 18040 10968 18068
rect 10827 18037 10839 18040
rect 10781 18031 10839 18037
rect 10962 18028 10968 18040
rect 11020 18028 11026 18080
rect 13354 18068 13360 18080
rect 13315 18040 13360 18068
rect 13354 18028 13360 18040
rect 13412 18028 13418 18080
rect 14458 18028 14464 18080
rect 14516 18068 14522 18080
rect 14645 18071 14703 18077
rect 14645 18068 14657 18071
rect 14516 18040 14657 18068
rect 14516 18028 14522 18040
rect 14645 18037 14657 18040
rect 14691 18037 14703 18071
rect 14645 18031 14703 18037
rect 18046 18028 18052 18080
rect 18104 18068 18110 18080
rect 19904 18068 19932 18108
rect 20530 18096 20536 18108
rect 20588 18096 20594 18148
rect 20622 18096 20628 18148
rect 20680 18136 20686 18148
rect 22646 18136 22652 18148
rect 20680 18108 22652 18136
rect 20680 18096 20686 18108
rect 22646 18096 22652 18108
rect 22704 18096 22710 18148
rect 18104 18040 19932 18068
rect 19981 18071 20039 18077
rect 18104 18028 18110 18040
rect 19981 18037 19993 18071
rect 20027 18068 20039 18071
rect 20438 18068 20444 18080
rect 20027 18040 20444 18068
rect 20027 18037 20039 18040
rect 19981 18031 20039 18037
rect 20438 18028 20444 18040
rect 20496 18028 20502 18080
rect 20714 18028 20720 18080
rect 20772 18068 20778 18080
rect 20901 18071 20959 18077
rect 20901 18068 20913 18071
rect 20772 18040 20913 18068
rect 20772 18028 20778 18040
rect 20901 18037 20913 18040
rect 20947 18037 20959 18071
rect 22848 18068 22876 18235
rect 23014 18232 23020 18235
rect 23072 18232 23078 18284
rect 23236 18281 23264 18312
rect 23477 18309 23489 18343
rect 23523 18340 23535 18343
rect 23998 18343 24056 18349
rect 23998 18340 24010 18343
rect 23523 18312 24010 18340
rect 23523 18309 23535 18312
rect 23477 18303 23535 18309
rect 23998 18309 24010 18312
rect 24044 18309 24056 18343
rect 23998 18303 24056 18309
rect 23109 18275 23167 18281
rect 23109 18241 23121 18275
rect 23155 18241 23167 18275
rect 23236 18275 23305 18281
rect 23236 18244 23259 18275
rect 23109 18235 23167 18241
rect 23247 18241 23259 18244
rect 23293 18241 23305 18275
rect 23247 18235 23305 18241
rect 23753 18275 23811 18281
rect 23753 18241 23765 18275
rect 23799 18272 23811 18275
rect 23842 18272 23848 18284
rect 23799 18244 23848 18272
rect 23799 18241 23811 18244
rect 23753 18235 23811 18241
rect 23124 18204 23152 18235
rect 23842 18232 23848 18244
rect 23900 18232 23906 18284
rect 23474 18204 23480 18216
rect 23124 18176 23480 18204
rect 23474 18164 23480 18176
rect 23532 18164 23538 18216
rect 22922 18068 22928 18080
rect 22848 18040 22928 18068
rect 20901 18031 20959 18037
rect 22922 18028 22928 18040
rect 22980 18028 22986 18080
rect 23106 18028 23112 18080
rect 23164 18068 23170 18080
rect 25133 18071 25191 18077
rect 25133 18068 25145 18071
rect 23164 18040 25145 18068
rect 23164 18028 23170 18040
rect 25133 18037 25145 18040
rect 25179 18037 25191 18071
rect 25133 18031 25191 18037
rect 1104 17978 28888 18000
rect 1104 17926 5582 17978
rect 5634 17926 5646 17978
rect 5698 17926 5710 17978
rect 5762 17926 5774 17978
rect 5826 17926 5838 17978
rect 5890 17926 14846 17978
rect 14898 17926 14910 17978
rect 14962 17926 14974 17978
rect 15026 17926 15038 17978
rect 15090 17926 15102 17978
rect 15154 17926 24110 17978
rect 24162 17926 24174 17978
rect 24226 17926 24238 17978
rect 24290 17926 24302 17978
rect 24354 17926 24366 17978
rect 24418 17926 28888 17978
rect 1104 17904 28888 17926
rect 8110 17864 8116 17876
rect 8071 17836 8116 17864
rect 8110 17824 8116 17836
rect 8168 17824 8174 17876
rect 10594 17864 10600 17876
rect 10555 17836 10600 17864
rect 10594 17824 10600 17836
rect 10652 17824 10658 17876
rect 11146 17864 11152 17876
rect 11107 17836 11152 17864
rect 11146 17824 11152 17836
rect 11204 17824 11210 17876
rect 12345 17867 12403 17873
rect 12345 17833 12357 17867
rect 12391 17864 12403 17867
rect 12710 17864 12716 17876
rect 12391 17836 12716 17864
rect 12391 17833 12403 17836
rect 12345 17827 12403 17833
rect 12710 17824 12716 17836
rect 12768 17864 12774 17876
rect 12805 17867 12863 17873
rect 12805 17864 12817 17867
rect 12768 17836 12817 17864
rect 12768 17824 12774 17836
rect 12805 17833 12817 17836
rect 12851 17864 12863 17867
rect 13354 17864 13360 17876
rect 12851 17836 13360 17864
rect 12851 17833 12863 17836
rect 12805 17827 12863 17833
rect 13354 17824 13360 17836
rect 13412 17864 13418 17876
rect 13449 17867 13507 17873
rect 13449 17864 13461 17867
rect 13412 17836 13461 17864
rect 13412 17824 13418 17836
rect 13449 17833 13461 17836
rect 13495 17833 13507 17867
rect 13449 17827 13507 17833
rect 17586 17824 17592 17876
rect 17644 17864 17650 17876
rect 17644 17836 18092 17864
rect 17644 17824 17650 17836
rect 10318 17796 10324 17808
rect 10231 17768 10324 17796
rect 10318 17756 10324 17768
rect 10376 17756 10382 17808
rect 12986 17796 12992 17808
rect 12947 17768 12992 17796
rect 12986 17756 12992 17768
rect 13044 17756 13050 17808
rect 13633 17799 13691 17805
rect 13633 17765 13645 17799
rect 13679 17796 13691 17799
rect 18064 17796 18092 17836
rect 18138 17824 18144 17876
rect 18196 17864 18202 17876
rect 18417 17867 18475 17873
rect 18417 17864 18429 17867
rect 18196 17836 18429 17864
rect 18196 17824 18202 17836
rect 18417 17833 18429 17836
rect 18463 17833 18475 17867
rect 18417 17827 18475 17833
rect 18598 17824 18604 17876
rect 18656 17864 18662 17876
rect 21177 17867 21235 17873
rect 21177 17864 21189 17867
rect 18656 17836 21189 17864
rect 18656 17824 18662 17836
rect 21177 17833 21189 17836
rect 21223 17864 21235 17867
rect 21634 17864 21640 17876
rect 21223 17836 21640 17864
rect 21223 17833 21235 17836
rect 21177 17827 21235 17833
rect 21634 17824 21640 17836
rect 21692 17824 21698 17876
rect 23014 17824 23020 17876
rect 23072 17864 23078 17876
rect 23293 17867 23351 17873
rect 23293 17864 23305 17867
rect 23072 17836 23305 17864
rect 23072 17824 23078 17836
rect 23293 17833 23305 17836
rect 23339 17833 23351 17867
rect 23293 17827 23351 17833
rect 13679 17768 15608 17796
rect 18064 17768 20484 17796
rect 13679 17765 13691 17768
rect 13633 17759 13691 17765
rect 10336 17728 10364 17756
rect 15470 17728 15476 17740
rect 10336 17700 13308 17728
rect 5994 17660 6000 17672
rect 5955 17632 6000 17660
rect 5994 17620 6000 17632
rect 6052 17620 6058 17672
rect 8941 17663 8999 17669
rect 8941 17629 8953 17663
rect 8987 17660 8999 17663
rect 9030 17660 9036 17672
rect 8987 17632 9036 17660
rect 8987 17629 8999 17632
rect 8941 17623 8999 17629
rect 9030 17620 9036 17632
rect 9088 17620 9094 17672
rect 10962 17660 10968 17672
rect 10923 17632 10968 17660
rect 10962 17620 10968 17632
rect 11020 17620 11026 17672
rect 11701 17663 11759 17669
rect 11701 17629 11713 17663
rect 11747 17660 11759 17663
rect 11974 17660 11980 17672
rect 11747 17632 11980 17660
rect 11747 17629 11759 17632
rect 11701 17623 11759 17629
rect 11974 17620 11980 17632
rect 12032 17620 12038 17672
rect 12161 17663 12219 17669
rect 12161 17629 12173 17663
rect 12207 17660 12219 17663
rect 12802 17660 12808 17672
rect 12207 17632 12808 17660
rect 12207 17629 12219 17632
rect 12161 17623 12219 17629
rect 12802 17620 12808 17632
rect 12860 17620 12866 17672
rect 6086 17552 6092 17604
rect 6144 17592 6150 17604
rect 6242 17595 6300 17601
rect 6242 17592 6254 17595
rect 6144 17564 6254 17592
rect 6144 17552 6150 17564
rect 6242 17561 6254 17564
rect 6288 17561 6300 17595
rect 8018 17592 8024 17604
rect 7979 17564 8024 17592
rect 6242 17555 6300 17561
rect 8018 17552 8024 17564
rect 8076 17552 8082 17604
rect 8662 17552 8668 17604
rect 8720 17592 8726 17604
rect 9186 17595 9244 17601
rect 9186 17592 9198 17595
rect 8720 17564 9198 17592
rect 8720 17552 8726 17564
rect 9186 17561 9198 17564
rect 9232 17561 9244 17595
rect 12618 17592 12624 17604
rect 12579 17564 12624 17592
rect 9186 17555 9244 17561
rect 12618 17552 12624 17564
rect 12676 17552 12682 17604
rect 13280 17601 13308 17700
rect 14568 17700 15148 17728
rect 15431 17700 15476 17728
rect 13495 17629 13553 17635
rect 13265 17595 13323 17601
rect 13265 17561 13277 17595
rect 13311 17561 13323 17595
rect 13495 17595 13507 17629
rect 13541 17604 13553 17629
rect 14182 17620 14188 17672
rect 14240 17660 14246 17672
rect 14323 17663 14381 17669
rect 14568 17666 14596 17700
rect 14323 17660 14335 17663
rect 14240 17632 14335 17660
rect 14240 17620 14246 17632
rect 14323 17629 14335 17632
rect 14369 17629 14381 17663
rect 14455 17654 14461 17666
rect 14323 17623 14381 17629
rect 14416 17626 14461 17654
rect 14455 17614 14461 17626
rect 14513 17614 14519 17666
rect 14553 17660 14611 17666
rect 14553 17626 14565 17660
rect 14599 17626 14611 17660
rect 14553 17620 14611 17626
rect 14642 17620 14648 17672
rect 14700 17660 14706 17672
rect 14737 17663 14795 17669
rect 14737 17660 14749 17663
rect 14700 17632 14749 17660
rect 14700 17620 14706 17632
rect 14737 17629 14749 17632
rect 14783 17660 14795 17663
rect 15013 17663 15071 17669
rect 15013 17660 15025 17663
rect 14783 17632 15025 17660
rect 14783 17629 14795 17632
rect 14737 17623 14795 17629
rect 15013 17629 15025 17632
rect 15059 17629 15071 17663
rect 15013 17623 15071 17629
rect 13541 17595 13544 17604
rect 13495 17592 13544 17595
rect 13265 17555 13323 17561
rect 13480 17564 13544 17592
rect 7374 17524 7380 17536
rect 7335 17496 7380 17524
rect 7374 17484 7380 17496
rect 7432 17484 7438 17536
rect 11885 17527 11943 17533
rect 11885 17493 11897 17527
rect 11931 17524 11943 17527
rect 12434 17524 12440 17536
rect 11931 17496 12440 17524
rect 11931 17493 11943 17496
rect 11885 17487 11943 17493
rect 12434 17484 12440 17496
rect 12492 17524 12498 17536
rect 12821 17527 12879 17533
rect 12821 17524 12833 17527
rect 12492 17496 12833 17524
rect 12492 17484 12498 17496
rect 12821 17493 12833 17496
rect 12867 17524 12879 17527
rect 13480 17524 13508 17564
rect 13538 17552 13544 17564
rect 13596 17552 13602 17604
rect 15120 17592 15148 17700
rect 15470 17688 15476 17700
rect 15528 17688 15534 17740
rect 15580 17728 15608 17768
rect 17957 17731 18015 17737
rect 15580 17700 15792 17728
rect 15194 17620 15200 17672
rect 15252 17660 15258 17672
rect 15381 17663 15439 17669
rect 15381 17660 15393 17663
rect 15252 17632 15393 17660
rect 15252 17620 15258 17632
rect 15381 17629 15393 17632
rect 15427 17629 15439 17663
rect 15654 17660 15660 17672
rect 15615 17632 15660 17660
rect 15381 17623 15439 17629
rect 15654 17620 15660 17632
rect 15712 17620 15718 17672
rect 15764 17669 15792 17700
rect 17957 17697 17969 17731
rect 18003 17728 18015 17731
rect 19334 17728 19340 17740
rect 18003 17700 19340 17728
rect 18003 17697 18015 17700
rect 17957 17691 18015 17697
rect 19334 17688 19340 17700
rect 19392 17688 19398 17740
rect 15749 17663 15807 17669
rect 15749 17629 15761 17663
rect 15795 17629 15807 17663
rect 19536 17660 19564 17768
rect 19797 17731 19855 17737
rect 19797 17697 19809 17731
rect 19843 17728 19855 17731
rect 19978 17728 19984 17740
rect 19843 17700 19984 17728
rect 19843 17697 19855 17700
rect 19797 17691 19855 17697
rect 19978 17688 19984 17700
rect 20036 17728 20042 17740
rect 20346 17728 20352 17740
rect 20036 17700 20352 17728
rect 20036 17688 20042 17700
rect 20346 17688 20352 17700
rect 20404 17688 20410 17740
rect 19613 17663 19671 17669
rect 19613 17660 19625 17663
rect 15749 17623 15807 17629
rect 15856 17632 19334 17660
rect 19536 17632 19625 17660
rect 15856 17592 15884 17632
rect 15120 17564 15884 17592
rect 15933 17595 15991 17601
rect 15933 17561 15945 17595
rect 15979 17592 15991 17595
rect 16482 17592 16488 17604
rect 15979 17564 16488 17592
rect 15979 17561 15991 17564
rect 15933 17555 15991 17561
rect 16482 17552 16488 17564
rect 16540 17552 16546 17604
rect 17712 17595 17770 17601
rect 17712 17561 17724 17595
rect 17758 17592 17770 17595
rect 18506 17592 18512 17604
rect 17758 17564 18512 17592
rect 17758 17561 17770 17564
rect 17712 17555 17770 17561
rect 18506 17552 18512 17564
rect 18564 17552 18570 17604
rect 18598 17552 18604 17604
rect 18656 17592 18662 17604
rect 18785 17595 18843 17601
rect 18656 17564 18701 17592
rect 18656 17552 18662 17564
rect 18785 17561 18797 17595
rect 18831 17561 18843 17595
rect 19306 17592 19334 17632
rect 19613 17629 19625 17632
rect 19659 17629 19671 17663
rect 19613 17623 19671 17629
rect 19705 17663 19763 17669
rect 19705 17629 19717 17663
rect 19751 17660 19763 17663
rect 19886 17660 19892 17672
rect 19751 17632 19892 17660
rect 19751 17629 19763 17632
rect 19705 17623 19763 17629
rect 19886 17620 19892 17632
rect 19944 17620 19950 17672
rect 20456 17657 20484 17768
rect 20622 17756 20628 17808
rect 20680 17756 20686 17808
rect 20714 17756 20720 17808
rect 20772 17756 20778 17808
rect 22278 17796 22284 17808
rect 22239 17768 22284 17796
rect 22278 17756 22284 17768
rect 22336 17756 22342 17808
rect 20637 17669 20665 17756
rect 20533 17663 20591 17669
rect 20533 17657 20545 17663
rect 20456 17629 20545 17657
rect 20579 17629 20591 17663
rect 20533 17623 20591 17629
rect 20622 17663 20680 17669
rect 20732 17666 20760 17756
rect 22738 17688 22744 17740
rect 22796 17728 22802 17740
rect 22796 17700 24532 17728
rect 22796 17688 22802 17700
rect 20622 17629 20634 17663
rect 20668 17629 20680 17663
rect 20622 17623 20680 17629
rect 20717 17660 20775 17666
rect 20717 17626 20729 17660
rect 20763 17626 20775 17660
rect 20717 17620 20775 17626
rect 20898 17620 20904 17672
rect 20956 17660 20962 17672
rect 21266 17660 21272 17672
rect 20956 17632 21272 17660
rect 20956 17620 20962 17632
rect 21266 17620 21272 17632
rect 21324 17620 21330 17672
rect 21821 17663 21879 17669
rect 21821 17629 21833 17663
rect 21867 17660 21879 17663
rect 23106 17660 23112 17672
rect 21867 17632 23112 17660
rect 21867 17629 21879 17632
rect 21821 17623 21879 17629
rect 23106 17620 23112 17632
rect 23164 17620 23170 17672
rect 19306 17564 20484 17592
rect 18785 17555 18843 17561
rect 14090 17524 14096 17536
rect 12867 17496 13508 17524
rect 14051 17496 14096 17524
rect 12867 17493 12879 17496
rect 12821 17487 12879 17493
rect 14090 17484 14096 17496
rect 14148 17484 14154 17536
rect 14642 17484 14648 17536
rect 14700 17524 14706 17536
rect 16114 17524 16120 17536
rect 14700 17496 16120 17524
rect 14700 17484 14706 17496
rect 16114 17484 16120 17496
rect 16172 17524 16178 17536
rect 16209 17527 16267 17533
rect 16209 17524 16221 17527
rect 16172 17496 16221 17524
rect 16172 17484 16178 17496
rect 16209 17493 16221 17496
rect 16255 17493 16267 17527
rect 16209 17487 16267 17493
rect 16298 17484 16304 17536
rect 16356 17524 16362 17536
rect 16577 17527 16635 17533
rect 16577 17524 16589 17527
rect 16356 17496 16589 17524
rect 16356 17484 16362 17496
rect 16577 17493 16589 17496
rect 16623 17524 16635 17527
rect 18230 17524 18236 17536
rect 16623 17496 18236 17524
rect 16623 17493 16635 17496
rect 16577 17487 16635 17493
rect 18230 17484 18236 17496
rect 18288 17484 18294 17536
rect 18800 17524 18828 17555
rect 19245 17527 19303 17533
rect 19245 17524 19257 17527
rect 18800 17496 19257 17524
rect 19245 17493 19257 17496
rect 19291 17493 19303 17527
rect 20254 17524 20260 17536
rect 20215 17496 20260 17524
rect 19245 17487 19303 17493
rect 20254 17484 20260 17496
rect 20312 17484 20318 17536
rect 20456 17524 20484 17564
rect 21726 17552 21732 17604
rect 21784 17592 21790 17604
rect 22005 17595 22063 17601
rect 22005 17592 22017 17595
rect 21784 17564 22017 17592
rect 21784 17552 21790 17564
rect 22005 17561 22017 17564
rect 22051 17561 22063 17595
rect 22462 17592 22468 17604
rect 22423 17564 22468 17592
rect 22005 17555 22063 17561
rect 22462 17552 22468 17564
rect 22520 17552 22526 17604
rect 22925 17595 22983 17601
rect 22925 17561 22937 17595
rect 22971 17561 22983 17595
rect 22925 17555 22983 17561
rect 21637 17527 21695 17533
rect 21637 17524 21649 17527
rect 20456 17496 21649 17524
rect 21637 17493 21649 17496
rect 21683 17493 21695 17527
rect 21637 17487 21695 17493
rect 21910 17484 21916 17536
rect 21968 17524 21974 17536
rect 22940 17524 22968 17555
rect 23014 17552 23020 17604
rect 23072 17592 23078 17604
rect 23753 17595 23811 17601
rect 23753 17592 23765 17595
rect 23072 17564 23765 17592
rect 23072 17552 23078 17564
rect 23753 17561 23765 17564
rect 23799 17561 23811 17595
rect 23753 17555 23811 17561
rect 23842 17552 23848 17604
rect 23900 17592 23906 17604
rect 23937 17595 23995 17601
rect 23937 17592 23949 17595
rect 23900 17564 23949 17592
rect 23900 17552 23906 17564
rect 23937 17561 23949 17564
rect 23983 17561 23995 17595
rect 23937 17555 23995 17561
rect 23198 17524 23204 17536
rect 21968 17496 23204 17524
rect 21968 17484 21974 17496
rect 23198 17484 23204 17496
rect 23256 17484 23262 17536
rect 23382 17484 23388 17536
rect 23440 17524 23446 17536
rect 24504 17533 24532 17700
rect 23569 17527 23627 17533
rect 23569 17524 23581 17527
rect 23440 17496 23581 17524
rect 23440 17484 23446 17496
rect 23569 17493 23581 17496
rect 23615 17493 23627 17527
rect 23569 17487 23627 17493
rect 24489 17527 24547 17533
rect 24489 17493 24501 17527
rect 24535 17524 24547 17527
rect 25406 17524 25412 17536
rect 24535 17496 25412 17524
rect 24535 17493 24547 17496
rect 24489 17487 24547 17493
rect 25406 17484 25412 17496
rect 25464 17484 25470 17536
rect 1104 17434 28888 17456
rect 1104 17382 10214 17434
rect 10266 17382 10278 17434
rect 10330 17382 10342 17434
rect 10394 17382 10406 17434
rect 10458 17382 10470 17434
rect 10522 17382 19478 17434
rect 19530 17382 19542 17434
rect 19594 17382 19606 17434
rect 19658 17382 19670 17434
rect 19722 17382 19734 17434
rect 19786 17382 28888 17434
rect 1104 17360 28888 17382
rect 5997 17323 6055 17329
rect 5997 17289 6009 17323
rect 6043 17320 6055 17323
rect 6086 17320 6092 17332
rect 6043 17292 6092 17320
rect 6043 17289 6055 17292
rect 5997 17283 6055 17289
rect 6086 17280 6092 17292
rect 6144 17280 6150 17332
rect 7009 17323 7067 17329
rect 7009 17320 7021 17323
rect 6886 17292 7021 17320
rect 5813 17187 5871 17193
rect 5813 17153 5825 17187
rect 5859 17184 5871 17187
rect 6365 17187 6423 17193
rect 6365 17184 6377 17187
rect 5859 17156 6377 17184
rect 5859 17153 5871 17156
rect 5813 17147 5871 17153
rect 6365 17153 6377 17156
rect 6411 17153 6423 17187
rect 6365 17147 6423 17153
rect 6549 17187 6607 17193
rect 6549 17153 6561 17187
rect 6595 17184 6607 17187
rect 6886 17184 6914 17292
rect 7009 17289 7021 17292
rect 7055 17289 7067 17323
rect 8662 17320 8668 17332
rect 8623 17292 8668 17320
rect 7009 17283 7067 17289
rect 8662 17280 8668 17292
rect 8720 17280 8726 17332
rect 9858 17320 9864 17332
rect 9819 17292 9864 17320
rect 9858 17280 9864 17292
rect 9916 17280 9922 17332
rect 13262 17320 13268 17332
rect 11348 17292 13268 17320
rect 7374 17252 7380 17264
rect 7287 17224 7380 17252
rect 7374 17212 7380 17224
rect 7432 17252 7438 17264
rect 9769 17255 9827 17261
rect 7432 17224 9444 17252
rect 7432 17212 7438 17224
rect 6595 17156 6914 17184
rect 8481 17187 8539 17193
rect 6595 17153 6607 17156
rect 6549 17147 6607 17153
rect 8481 17153 8493 17187
rect 8527 17184 8539 17187
rect 8941 17187 8999 17193
rect 8941 17184 8953 17187
rect 8527 17156 8953 17184
rect 8527 17153 8539 17156
rect 8481 17147 8539 17153
rect 8941 17153 8953 17156
rect 8987 17153 8999 17187
rect 9122 17184 9128 17196
rect 9083 17156 9128 17184
rect 8941 17147 8999 17153
rect 9122 17144 9128 17156
rect 9180 17144 9186 17196
rect 6638 17076 6644 17128
rect 6696 17116 6702 17128
rect 6733 17119 6791 17125
rect 6733 17116 6745 17119
rect 6696 17088 6745 17116
rect 6696 17076 6702 17088
rect 6733 17085 6745 17088
rect 6779 17085 6791 17119
rect 7466 17116 7472 17128
rect 7427 17088 7472 17116
rect 6733 17079 6791 17085
rect 7466 17076 7472 17088
rect 7524 17076 7530 17128
rect 7653 17119 7711 17125
rect 7653 17085 7665 17119
rect 7699 17116 7711 17119
rect 7834 17116 7840 17128
rect 7699 17088 7840 17116
rect 7699 17085 7711 17088
rect 7653 17079 7711 17085
rect 7834 17076 7840 17088
rect 7892 17116 7898 17128
rect 8018 17116 8024 17128
rect 7892 17088 8024 17116
rect 7892 17076 7898 17088
rect 8018 17076 8024 17088
rect 8076 17076 8082 17128
rect 9306 17116 9312 17128
rect 9267 17088 9312 17116
rect 9306 17076 9312 17088
rect 9364 17076 9370 17128
rect 9416 17116 9444 17224
rect 9769 17221 9781 17255
rect 9815 17252 9827 17255
rect 10594 17252 10600 17264
rect 9815 17224 10600 17252
rect 9815 17221 9827 17224
rect 9769 17215 9827 17221
rect 10594 17212 10600 17224
rect 10652 17252 10658 17264
rect 10962 17252 10968 17264
rect 10652 17224 10968 17252
rect 10652 17212 10658 17224
rect 10962 17212 10968 17224
rect 11020 17212 11026 17264
rect 10689 17187 10747 17193
rect 10689 17153 10701 17187
rect 10735 17184 10747 17187
rect 11348 17184 11376 17292
rect 13262 17280 13268 17292
rect 13320 17280 13326 17332
rect 14737 17323 14795 17329
rect 14737 17289 14749 17323
rect 14783 17320 14795 17323
rect 15562 17320 15568 17332
rect 14783 17292 15568 17320
rect 14783 17289 14795 17292
rect 14737 17283 14795 17289
rect 15562 17280 15568 17292
rect 15620 17280 15626 17332
rect 17497 17323 17555 17329
rect 17497 17289 17509 17323
rect 17543 17320 17555 17323
rect 18230 17320 18236 17332
rect 17543 17292 18236 17320
rect 17543 17289 17555 17292
rect 17497 17283 17555 17289
rect 18230 17280 18236 17292
rect 18288 17280 18294 17332
rect 18506 17280 18512 17332
rect 18564 17320 18570 17332
rect 18693 17323 18751 17329
rect 18693 17320 18705 17323
rect 18564 17292 18705 17320
rect 18564 17280 18570 17292
rect 18693 17289 18705 17292
rect 18739 17289 18751 17323
rect 18693 17283 18751 17289
rect 20993 17323 21051 17329
rect 20993 17289 21005 17323
rect 21039 17320 21051 17323
rect 21082 17320 21088 17332
rect 21039 17292 21088 17320
rect 21039 17289 21051 17292
rect 20993 17283 21051 17289
rect 21082 17280 21088 17292
rect 21140 17280 21146 17332
rect 23014 17280 23020 17332
rect 23072 17320 23078 17332
rect 25317 17323 25375 17329
rect 25317 17320 25329 17323
rect 23072 17292 25329 17320
rect 23072 17280 23078 17292
rect 25317 17289 25329 17292
rect 25363 17289 25375 17323
rect 25317 17283 25375 17289
rect 25406 17280 25412 17332
rect 25464 17320 25470 17332
rect 28169 17323 28227 17329
rect 28169 17320 28181 17323
rect 25464 17292 28181 17320
rect 25464 17280 25470 17292
rect 28169 17289 28181 17292
rect 28215 17289 28227 17323
rect 28169 17283 28227 17289
rect 11606 17212 11612 17264
rect 11664 17252 11670 17264
rect 11762 17255 11820 17261
rect 11762 17252 11774 17255
rect 11664 17224 11774 17252
rect 11664 17212 11670 17224
rect 11762 17221 11774 17224
rect 11808 17221 11820 17255
rect 11762 17215 11820 17221
rect 12342 17212 12348 17264
rect 12400 17252 12406 17264
rect 13173 17255 13231 17261
rect 13173 17252 13185 17255
rect 12400 17224 13185 17252
rect 12400 17212 12406 17224
rect 13173 17221 13185 17224
rect 13219 17221 13231 17255
rect 13173 17215 13231 17221
rect 13357 17255 13415 17261
rect 13357 17221 13369 17255
rect 13403 17252 13415 17255
rect 14921 17255 14979 17261
rect 14921 17252 14933 17255
rect 13403 17224 14933 17252
rect 13403 17221 13415 17224
rect 13357 17215 13415 17221
rect 14921 17221 14933 17224
rect 14967 17221 14979 17255
rect 14921 17215 14979 17221
rect 15105 17255 15163 17261
rect 15105 17221 15117 17255
rect 15151 17252 15163 17255
rect 16945 17255 17003 17261
rect 15151 17224 16068 17252
rect 15151 17221 15163 17224
rect 15105 17215 15163 17221
rect 10735 17156 11376 17184
rect 10735 17153 10747 17156
rect 10689 17147 10747 17153
rect 12250 17144 12256 17196
rect 12308 17184 12314 17196
rect 13372 17184 13400 17215
rect 12308 17156 13400 17184
rect 12308 17144 12314 17156
rect 13998 17144 14004 17196
rect 14056 17184 14062 17196
rect 14093 17187 14151 17193
rect 14093 17184 14105 17187
rect 14056 17156 14105 17184
rect 14056 17144 14062 17156
rect 14093 17153 14105 17156
rect 14139 17153 14151 17187
rect 14093 17147 14151 17153
rect 14185 17187 14243 17193
rect 14185 17153 14197 17187
rect 14231 17153 14243 17187
rect 14185 17147 14243 17153
rect 14277 17187 14335 17193
rect 14277 17153 14289 17187
rect 14323 17153 14335 17187
rect 14458 17184 14464 17196
rect 14419 17156 14464 17184
rect 14277 17147 14335 17153
rect 10781 17119 10839 17125
rect 10781 17116 10793 17119
rect 9416 17088 10793 17116
rect 10781 17085 10793 17088
rect 10827 17085 10839 17119
rect 10781 17079 10839 17085
rect 10965 17119 11023 17125
rect 10965 17085 10977 17119
rect 11011 17116 11023 17119
rect 11054 17116 11060 17128
rect 11011 17088 11060 17116
rect 11011 17085 11023 17088
rect 10965 17079 11023 17085
rect 11054 17076 11060 17088
rect 11112 17076 11118 17128
rect 11514 17116 11520 17128
rect 11427 17088 11520 17116
rect 11514 17076 11520 17088
rect 11572 17076 11578 17128
rect 13630 17076 13636 17128
rect 13688 17116 13694 17128
rect 14200 17116 14228 17147
rect 13688 17088 14228 17116
rect 13688 17076 13694 17088
rect 1394 17048 1400 17060
rect 1355 17020 1400 17048
rect 1394 17008 1400 17020
rect 1452 17008 1458 17060
rect 10318 16980 10324 16992
rect 10279 16952 10324 16980
rect 10318 16940 10324 16952
rect 10376 16940 10382 16992
rect 11532 16980 11560 17076
rect 12986 17008 12992 17060
rect 13044 17048 13050 17060
rect 14292 17048 14320 17147
rect 14458 17144 14464 17156
rect 14516 17144 14522 17196
rect 15381 17187 15439 17193
rect 15381 17153 15393 17187
rect 15427 17184 15439 17187
rect 15746 17184 15752 17196
rect 15427 17156 15752 17184
rect 15427 17153 15439 17156
rect 15381 17147 15439 17153
rect 15746 17144 15752 17156
rect 15804 17144 15810 17196
rect 14550 17076 14556 17128
rect 14608 17116 14614 17128
rect 15470 17116 15476 17128
rect 14608 17088 15476 17116
rect 14608 17076 14614 17088
rect 15470 17076 15476 17088
rect 15528 17116 15534 17128
rect 15657 17119 15715 17125
rect 15657 17116 15669 17119
rect 15528 17088 15669 17116
rect 15528 17076 15534 17088
rect 15657 17085 15669 17088
rect 15703 17085 15715 17119
rect 16040 17116 16068 17224
rect 16945 17221 16957 17255
rect 16991 17252 17003 17255
rect 19880 17255 19938 17261
rect 16991 17224 18552 17252
rect 16991 17221 17003 17224
rect 16945 17215 17003 17221
rect 16114 17144 16120 17196
rect 16172 17184 16178 17196
rect 17586 17184 17592 17196
rect 16172 17156 17448 17184
rect 17547 17156 17592 17184
rect 16172 17144 16178 17156
rect 17218 17116 17224 17128
rect 16040 17088 17224 17116
rect 15657 17079 15715 17085
rect 17218 17076 17224 17088
rect 17276 17116 17282 17128
rect 17313 17119 17371 17125
rect 17313 17116 17325 17119
rect 17276 17088 17325 17116
rect 17276 17076 17282 17088
rect 17313 17085 17325 17088
rect 17359 17085 17371 17119
rect 17420 17116 17448 17156
rect 17586 17144 17592 17156
rect 17644 17144 17650 17196
rect 17954 17144 17960 17196
rect 18012 17184 18018 17196
rect 18524 17193 18552 17224
rect 19880 17221 19892 17255
rect 19926 17252 19938 17255
rect 20254 17252 20260 17264
rect 19926 17224 20260 17252
rect 19926 17221 19938 17224
rect 19880 17215 19938 17221
rect 20254 17212 20260 17224
rect 20312 17212 20318 17264
rect 21468 17224 22232 17252
rect 18233 17187 18291 17193
rect 18233 17184 18245 17187
rect 18012 17156 18245 17184
rect 18012 17144 18018 17156
rect 18233 17153 18245 17156
rect 18279 17153 18291 17187
rect 18233 17147 18291 17153
rect 18509 17187 18567 17193
rect 18509 17153 18521 17187
rect 18555 17184 18567 17187
rect 18690 17184 18696 17196
rect 18555 17156 18696 17184
rect 18555 17153 18567 17156
rect 18509 17147 18567 17153
rect 18690 17144 18696 17156
rect 18748 17144 18754 17196
rect 19334 17144 19340 17196
rect 19392 17184 19398 17196
rect 19613 17187 19671 17193
rect 19613 17184 19625 17187
rect 19392 17156 19625 17184
rect 19392 17144 19398 17156
rect 19613 17153 19625 17156
rect 19659 17153 19671 17187
rect 21174 17184 21180 17196
rect 19613 17147 19671 17153
rect 19720 17156 21180 17184
rect 19720 17116 19748 17156
rect 21174 17144 21180 17156
rect 21232 17184 21238 17196
rect 21358 17184 21364 17196
rect 21232 17156 21364 17184
rect 21232 17144 21238 17156
rect 21358 17144 21364 17156
rect 21416 17144 21422 17196
rect 21468 17193 21496 17224
rect 22204 17196 22232 17224
rect 21453 17187 21511 17193
rect 21453 17153 21465 17187
rect 21499 17153 21511 17187
rect 21453 17147 21511 17153
rect 22005 17187 22063 17193
rect 22005 17153 22017 17187
rect 22051 17153 22063 17187
rect 22186 17184 22192 17196
rect 22147 17156 22192 17184
rect 22005 17147 22063 17153
rect 17420 17088 19748 17116
rect 22020 17116 22048 17147
rect 22186 17144 22192 17156
rect 22244 17144 22250 17196
rect 23198 17184 23204 17196
rect 23159 17156 23204 17184
rect 23198 17144 23204 17156
rect 23256 17144 23262 17196
rect 23842 17144 23848 17196
rect 23900 17184 23906 17196
rect 24193 17187 24251 17193
rect 24193 17184 24205 17187
rect 23900 17156 24205 17184
rect 23900 17144 23906 17156
rect 24193 17153 24205 17156
rect 24239 17153 24251 17187
rect 24193 17147 24251 17153
rect 27801 17187 27859 17193
rect 27801 17153 27813 17187
rect 27847 17184 27859 17187
rect 28350 17184 28356 17196
rect 27847 17156 28356 17184
rect 27847 17153 27859 17156
rect 27801 17147 27859 17153
rect 28350 17144 28356 17156
rect 28408 17144 28414 17196
rect 23014 17116 23020 17128
rect 22020 17088 23020 17116
rect 17313 17079 17371 17085
rect 23014 17076 23020 17088
rect 23072 17076 23078 17128
rect 23477 17119 23535 17125
rect 23477 17085 23489 17119
rect 23523 17116 23535 17119
rect 23750 17116 23756 17128
rect 23523 17088 23756 17116
rect 23523 17085 23535 17088
rect 23477 17079 23535 17085
rect 23750 17076 23756 17088
rect 23808 17076 23814 17128
rect 23934 17116 23940 17128
rect 23895 17088 23940 17116
rect 23934 17076 23940 17088
rect 23992 17076 23998 17128
rect 19610 17048 19616 17060
rect 13044 17020 14136 17048
rect 14292 17020 19616 17048
rect 13044 17008 13050 17020
rect 11882 16980 11888 16992
rect 11532 16952 11888 16980
rect 11882 16940 11888 16952
rect 11940 16940 11946 16992
rect 12897 16983 12955 16989
rect 12897 16949 12909 16983
rect 12943 16980 12955 16983
rect 13262 16980 13268 16992
rect 12943 16952 13268 16980
rect 12943 16949 12955 16952
rect 12897 16943 12955 16949
rect 13262 16940 13268 16952
rect 13320 16940 13326 16992
rect 13814 16980 13820 16992
rect 13775 16952 13820 16980
rect 13814 16940 13820 16952
rect 13872 16940 13878 16992
rect 14108 16980 14136 17020
rect 19610 17008 19616 17020
rect 19668 17008 19674 17060
rect 14458 16980 14464 16992
rect 14108 16952 14464 16980
rect 14458 16940 14464 16952
rect 14516 16940 14522 16992
rect 15194 16940 15200 16992
rect 15252 16980 15258 16992
rect 17494 16980 17500 16992
rect 15252 16952 17500 16980
rect 15252 16940 15258 16952
rect 17494 16940 17500 16952
rect 17552 16940 17558 16992
rect 17957 16983 18015 16989
rect 17957 16949 17969 16983
rect 18003 16980 18015 16983
rect 18325 16983 18383 16989
rect 18325 16980 18337 16983
rect 18003 16952 18337 16980
rect 18003 16949 18015 16952
rect 17957 16943 18015 16949
rect 18325 16949 18337 16952
rect 18371 16949 18383 16983
rect 19058 16980 19064 16992
rect 19019 16952 19064 16980
rect 18325 16943 18383 16949
rect 19058 16940 19064 16952
rect 19116 16940 19122 16992
rect 19518 16940 19524 16992
rect 19576 16980 19582 16992
rect 20346 16980 20352 16992
rect 19576 16952 20352 16980
rect 19576 16940 19582 16952
rect 20346 16940 20352 16952
rect 20404 16940 20410 16992
rect 20714 16940 20720 16992
rect 20772 16980 20778 16992
rect 21269 16983 21327 16989
rect 21269 16980 21281 16983
rect 20772 16952 21281 16980
rect 20772 16940 20778 16952
rect 21269 16949 21281 16952
rect 21315 16980 21327 16983
rect 21726 16980 21732 16992
rect 21315 16952 21732 16980
rect 21315 16949 21327 16952
rect 21269 16943 21327 16949
rect 21726 16940 21732 16952
rect 21784 16940 21790 16992
rect 21821 16983 21879 16989
rect 21821 16949 21833 16983
rect 21867 16980 21879 16983
rect 21910 16980 21916 16992
rect 21867 16952 21916 16980
rect 21867 16949 21879 16952
rect 21821 16943 21879 16949
rect 21910 16940 21916 16952
rect 21968 16940 21974 16992
rect 1104 16890 28888 16912
rect 1104 16838 5582 16890
rect 5634 16838 5646 16890
rect 5698 16838 5710 16890
rect 5762 16838 5774 16890
rect 5826 16838 5838 16890
rect 5890 16838 14846 16890
rect 14898 16838 14910 16890
rect 14962 16838 14974 16890
rect 15026 16838 15038 16890
rect 15090 16838 15102 16890
rect 15154 16838 24110 16890
rect 24162 16838 24174 16890
rect 24226 16838 24238 16890
rect 24290 16838 24302 16890
rect 24354 16838 24366 16890
rect 24418 16838 28888 16890
rect 1104 16816 28888 16838
rect 7193 16779 7251 16785
rect 7193 16745 7205 16779
rect 7239 16776 7251 16779
rect 7466 16776 7472 16788
rect 7239 16748 7472 16776
rect 7239 16745 7251 16748
rect 7193 16739 7251 16745
rect 7466 16736 7472 16748
rect 7524 16776 7530 16788
rect 7650 16776 7656 16788
rect 7524 16748 7656 16776
rect 7524 16736 7530 16748
rect 7650 16736 7656 16748
rect 7708 16776 7714 16788
rect 7708 16748 9168 16776
rect 7708 16736 7714 16748
rect 8573 16643 8631 16649
rect 8573 16609 8585 16643
rect 8619 16640 8631 16643
rect 9030 16640 9036 16652
rect 8619 16612 9036 16640
rect 8619 16609 8631 16612
rect 8573 16603 8631 16609
rect 9030 16600 9036 16612
rect 9088 16600 9094 16652
rect 9140 16640 9168 16748
rect 9858 16736 9864 16788
rect 9916 16776 9922 16788
rect 10686 16776 10692 16788
rect 9916 16748 10692 16776
rect 9916 16736 9922 16748
rect 10686 16736 10692 16748
rect 10744 16736 10750 16788
rect 10781 16779 10839 16785
rect 10781 16745 10793 16779
rect 10827 16776 10839 16779
rect 10870 16776 10876 16788
rect 10827 16748 10876 16776
rect 10827 16745 10839 16748
rect 10781 16739 10839 16745
rect 10870 16736 10876 16748
rect 10928 16736 10934 16788
rect 11054 16736 11060 16788
rect 11112 16776 11118 16788
rect 11149 16779 11207 16785
rect 11149 16776 11161 16779
rect 11112 16748 11161 16776
rect 11112 16736 11118 16748
rect 11149 16745 11161 16748
rect 11195 16745 11207 16779
rect 12158 16776 12164 16788
rect 12119 16748 12164 16776
rect 11149 16739 11207 16745
rect 12158 16736 12164 16748
rect 12216 16776 12222 16788
rect 15838 16776 15844 16788
rect 12216 16748 15844 16776
rect 12216 16736 12222 16748
rect 15838 16736 15844 16748
rect 15896 16736 15902 16788
rect 16850 16776 16856 16788
rect 16811 16748 16856 16776
rect 16850 16736 16856 16748
rect 16908 16736 16914 16788
rect 17218 16776 17224 16788
rect 17179 16748 17224 16776
rect 17218 16736 17224 16748
rect 17276 16736 17282 16788
rect 18322 16736 18328 16788
rect 18380 16776 18386 16788
rect 19242 16776 19248 16788
rect 18380 16748 19248 16776
rect 18380 16736 18386 16748
rect 19242 16736 19248 16748
rect 19300 16736 19306 16788
rect 19518 16776 19524 16788
rect 19479 16748 19524 16776
rect 19518 16736 19524 16748
rect 19576 16736 19582 16788
rect 19610 16736 19616 16788
rect 19668 16776 19674 16788
rect 20349 16779 20407 16785
rect 20349 16776 20361 16779
rect 19668 16748 20361 16776
rect 19668 16736 19674 16748
rect 20349 16745 20361 16748
rect 20395 16745 20407 16779
rect 23842 16776 23848 16788
rect 23803 16748 23848 16776
rect 20349 16739 20407 16745
rect 23842 16736 23848 16748
rect 23900 16736 23906 16788
rect 25038 16776 25044 16788
rect 24999 16748 25044 16776
rect 25038 16736 25044 16748
rect 25096 16736 25102 16788
rect 11072 16708 11100 16736
rect 9876 16680 11100 16708
rect 9876 16649 9904 16680
rect 13630 16668 13636 16720
rect 13688 16708 13694 16720
rect 14093 16711 14151 16717
rect 14093 16708 14105 16711
rect 13688 16680 14105 16708
rect 13688 16668 13694 16680
rect 14093 16677 14105 16680
rect 14139 16677 14151 16711
rect 14921 16711 14979 16717
rect 14921 16708 14933 16711
rect 14093 16671 14151 16677
rect 14292 16680 14933 16708
rect 9677 16643 9735 16649
rect 9677 16640 9689 16643
rect 9140 16612 9689 16640
rect 9677 16609 9689 16612
rect 9723 16609 9735 16643
rect 9677 16603 9735 16609
rect 9861 16643 9919 16649
rect 9861 16609 9873 16643
rect 9907 16609 9919 16643
rect 9861 16603 9919 16609
rect 10318 16600 10324 16652
rect 10376 16640 10382 16652
rect 12529 16643 12587 16649
rect 10376 16612 10640 16640
rect 10376 16600 10382 16612
rect 1673 16575 1731 16581
rect 1673 16541 1685 16575
rect 1719 16572 1731 16575
rect 4614 16572 4620 16584
rect 1719 16544 4620 16572
rect 1719 16541 1731 16544
rect 1673 16535 1731 16541
rect 4614 16532 4620 16544
rect 4672 16532 4678 16584
rect 9306 16532 9312 16584
rect 9364 16572 9370 16584
rect 9766 16572 9772 16584
rect 9364 16544 9772 16572
rect 9364 16532 9370 16544
rect 9766 16532 9772 16544
rect 9824 16572 9830 16584
rect 10612 16581 10640 16612
rect 12529 16609 12541 16643
rect 12575 16640 12587 16643
rect 13906 16640 13912 16652
rect 12575 16612 13912 16640
rect 12575 16609 12587 16612
rect 12529 16603 12587 16609
rect 13906 16600 13912 16612
rect 13964 16600 13970 16652
rect 10505 16575 10563 16581
rect 10505 16572 10517 16575
rect 9824 16544 10517 16572
rect 9824 16532 9830 16544
rect 10505 16541 10517 16544
rect 10551 16541 10563 16575
rect 10505 16535 10563 16541
rect 10597 16575 10655 16581
rect 10597 16541 10609 16575
rect 10643 16574 10655 16575
rect 10643 16546 10677 16574
rect 10643 16541 10655 16546
rect 10597 16535 10655 16541
rect 8294 16504 8300 16516
rect 8352 16513 8358 16516
rect 8264 16476 8300 16504
rect 8294 16464 8300 16476
rect 8352 16467 8364 16513
rect 10520 16504 10548 16535
rect 10778 16532 10784 16584
rect 10836 16572 10842 16584
rect 11701 16575 11759 16581
rect 11701 16572 11713 16575
rect 10836 16544 11713 16572
rect 10836 16532 10842 16544
rect 11701 16541 11713 16544
rect 11747 16541 11759 16575
rect 11701 16535 11759 16541
rect 12713 16575 12771 16581
rect 12713 16541 12725 16575
rect 12759 16541 12771 16575
rect 12713 16535 12771 16541
rect 12989 16575 13047 16581
rect 12989 16541 13001 16575
rect 13035 16572 13047 16575
rect 13265 16575 13323 16581
rect 13265 16572 13277 16575
rect 13035 16544 13277 16572
rect 13035 16541 13047 16544
rect 12989 16535 13047 16541
rect 13265 16541 13277 16544
rect 13311 16541 13323 16575
rect 13265 16535 13323 16541
rect 10870 16504 10876 16516
rect 10520 16476 10876 16504
rect 8352 16464 8358 16467
rect 10870 16464 10876 16476
rect 10928 16464 10934 16516
rect 11146 16464 11152 16516
rect 11204 16504 11210 16516
rect 11241 16507 11299 16513
rect 11241 16504 11253 16507
rect 11204 16476 11253 16504
rect 11204 16464 11210 16476
rect 11241 16473 11253 16476
rect 11287 16473 11299 16507
rect 11882 16504 11888 16516
rect 11843 16476 11888 16504
rect 11241 16467 11299 16473
rect 11882 16464 11888 16476
rect 11940 16464 11946 16516
rect 12728 16504 12756 16535
rect 13280 16504 13308 16535
rect 13354 16532 13360 16584
rect 13412 16572 13418 16584
rect 13412 16544 13457 16572
rect 13412 16532 13418 16544
rect 13538 16532 13544 16584
rect 13596 16572 13602 16584
rect 14090 16572 14096 16584
rect 13596 16544 14096 16572
rect 13596 16532 13602 16544
rect 14090 16532 14096 16544
rect 14148 16532 14154 16584
rect 14292 16581 14320 16680
rect 14921 16677 14933 16680
rect 14967 16677 14979 16711
rect 14921 16671 14979 16677
rect 15010 16668 15016 16720
rect 15068 16708 15074 16720
rect 16209 16711 16267 16717
rect 15068 16680 16068 16708
rect 15068 16668 15074 16680
rect 14550 16640 14556 16652
rect 14511 16612 14556 16640
rect 14550 16600 14556 16612
rect 14608 16600 14614 16652
rect 15746 16640 15752 16652
rect 15707 16612 15752 16640
rect 15746 16600 15752 16612
rect 15804 16600 15810 16652
rect 14277 16575 14335 16581
rect 14277 16541 14289 16575
rect 14323 16541 14335 16575
rect 14277 16535 14335 16541
rect 14366 16532 14372 16584
rect 14424 16572 14430 16584
rect 14642 16572 14648 16584
rect 14424 16544 14469 16572
rect 14603 16544 14648 16572
rect 14424 16532 14430 16544
rect 14642 16532 14648 16544
rect 14700 16532 14706 16584
rect 15102 16572 15108 16584
rect 15063 16544 15108 16572
rect 15102 16532 15108 16544
rect 15160 16532 15166 16584
rect 15381 16575 15439 16581
rect 15381 16572 15393 16575
rect 15212 16544 15393 16572
rect 15212 16504 15240 16544
rect 15381 16541 15393 16544
rect 15427 16572 15439 16575
rect 15470 16572 15476 16584
rect 15427 16544 15476 16572
rect 15427 16541 15439 16544
rect 15381 16535 15439 16541
rect 15470 16532 15476 16544
rect 15528 16532 15534 16584
rect 15654 16572 15660 16584
rect 15615 16544 15660 16572
rect 15654 16532 15660 16544
rect 15712 16532 15718 16584
rect 15930 16572 15936 16584
rect 15891 16544 15936 16572
rect 15930 16532 15936 16544
rect 15988 16532 15994 16584
rect 16040 16581 16068 16680
rect 16209 16677 16221 16711
rect 16255 16708 16267 16711
rect 22646 16708 22652 16720
rect 16255 16680 21956 16708
rect 22607 16680 22652 16708
rect 16255 16677 16267 16680
rect 16209 16671 16267 16677
rect 16945 16643 17003 16649
rect 16945 16609 16957 16643
rect 16991 16640 17003 16643
rect 17310 16640 17316 16652
rect 16991 16612 17316 16640
rect 16991 16609 17003 16612
rect 16945 16603 17003 16609
rect 17310 16600 17316 16612
rect 17368 16600 17374 16652
rect 18141 16643 18199 16649
rect 18141 16640 18153 16643
rect 17420 16612 18153 16640
rect 16025 16575 16083 16581
rect 16025 16541 16037 16575
rect 16071 16541 16083 16575
rect 16025 16535 16083 16541
rect 17037 16575 17095 16581
rect 17037 16541 17049 16575
rect 17083 16541 17095 16575
rect 17037 16535 17095 16541
rect 12728 16476 13032 16504
rect 13280 16476 15240 16504
rect 15289 16507 15347 16513
rect 1486 16436 1492 16448
rect 1447 16408 1492 16436
rect 1486 16396 1492 16408
rect 1544 16396 1550 16448
rect 9214 16436 9220 16448
rect 9175 16408 9220 16436
rect 9214 16396 9220 16408
rect 9272 16396 9278 16448
rect 9585 16439 9643 16445
rect 9585 16405 9597 16439
rect 9631 16436 9643 16439
rect 10686 16436 10692 16448
rect 9631 16408 10692 16436
rect 9631 16405 9643 16408
rect 9585 16399 9643 16405
rect 10686 16396 10692 16408
rect 10744 16396 10750 16448
rect 12894 16436 12900 16448
rect 12855 16408 12900 16436
rect 12894 16396 12900 16408
rect 12952 16396 12958 16448
rect 13004 16436 13032 16476
rect 15289 16473 15301 16507
rect 15335 16504 15347 16507
rect 16298 16504 16304 16516
rect 15335 16476 16304 16504
rect 15335 16473 15347 16476
rect 15289 16467 15347 16473
rect 16298 16464 16304 16476
rect 16356 16464 16362 16516
rect 16758 16504 16764 16516
rect 16719 16476 16764 16504
rect 16758 16464 16764 16476
rect 16816 16464 16822 16516
rect 17052 16504 17080 16535
rect 17218 16532 17224 16584
rect 17276 16572 17282 16584
rect 17420 16572 17448 16612
rect 18141 16609 18153 16612
rect 18187 16609 18199 16643
rect 20254 16640 20260 16652
rect 18141 16603 18199 16609
rect 18248 16612 20260 16640
rect 17276 16544 17448 16572
rect 18049 16575 18107 16581
rect 17276 16532 17282 16544
rect 18049 16541 18061 16575
rect 18095 16572 18107 16575
rect 18248 16572 18276 16612
rect 20254 16600 20260 16612
rect 20312 16600 20318 16652
rect 21928 16640 21956 16680
rect 22646 16668 22652 16680
rect 22704 16668 22710 16720
rect 21928 16612 22048 16640
rect 18095 16544 18276 16572
rect 18601 16575 18659 16581
rect 18095 16541 18107 16544
rect 18049 16535 18107 16541
rect 18601 16541 18613 16575
rect 18647 16572 18659 16575
rect 19242 16572 19248 16584
rect 18647 16544 18920 16572
rect 19203 16544 19248 16572
rect 18647 16541 18659 16544
rect 18601 16535 18659 16541
rect 18414 16504 18420 16516
rect 17052 16476 18420 16504
rect 18414 16464 18420 16476
rect 18472 16464 18478 16516
rect 13538 16436 13544 16448
rect 13004 16408 13544 16436
rect 13538 16396 13544 16408
rect 13596 16396 13602 16448
rect 13725 16439 13783 16445
rect 13725 16405 13737 16439
rect 13771 16436 13783 16439
rect 15102 16436 15108 16448
rect 13771 16408 15108 16436
rect 13771 16405 13783 16408
rect 13725 16399 13783 16405
rect 15102 16396 15108 16408
rect 15160 16396 15166 16448
rect 15194 16396 15200 16448
rect 15252 16436 15258 16448
rect 16390 16436 16396 16448
rect 15252 16408 16396 16436
rect 15252 16396 15258 16408
rect 16390 16396 16396 16408
rect 16448 16396 16454 16448
rect 17589 16439 17647 16445
rect 17589 16405 17601 16439
rect 17635 16436 17647 16439
rect 17770 16436 17776 16448
rect 17635 16408 17776 16436
rect 17635 16405 17647 16408
rect 17589 16399 17647 16405
rect 17770 16396 17776 16408
rect 17828 16396 17834 16448
rect 17957 16439 18015 16445
rect 17957 16405 17969 16439
rect 18003 16436 18015 16439
rect 18046 16436 18052 16448
rect 18003 16408 18052 16436
rect 18003 16405 18015 16408
rect 17957 16399 18015 16405
rect 18046 16396 18052 16408
rect 18104 16436 18110 16448
rect 18230 16436 18236 16448
rect 18104 16408 18236 16436
rect 18104 16396 18110 16408
rect 18230 16396 18236 16408
rect 18288 16396 18294 16448
rect 18690 16396 18696 16448
rect 18748 16436 18754 16448
rect 18785 16439 18843 16445
rect 18785 16436 18797 16439
rect 18748 16408 18797 16436
rect 18748 16396 18754 16408
rect 18785 16405 18797 16408
rect 18831 16405 18843 16439
rect 18892 16436 18920 16544
rect 19242 16532 19248 16544
rect 19300 16532 19306 16584
rect 19521 16575 19579 16581
rect 19521 16541 19533 16575
rect 19567 16541 19579 16575
rect 20162 16572 20168 16584
rect 19521 16535 19579 16541
rect 19628 16544 20168 16572
rect 19058 16464 19064 16516
rect 19116 16504 19122 16516
rect 19536 16504 19564 16535
rect 19116 16476 19564 16504
rect 19116 16464 19122 16476
rect 19628 16436 19656 16544
rect 20162 16532 20168 16544
rect 20220 16532 20226 16584
rect 20533 16575 20591 16581
rect 20533 16541 20545 16575
rect 20579 16572 20591 16575
rect 21082 16572 21088 16584
rect 20579 16544 21088 16572
rect 20579 16541 20591 16544
rect 20533 16535 20591 16541
rect 21082 16532 21088 16544
rect 21140 16532 21146 16584
rect 21726 16572 21732 16584
rect 21687 16544 21732 16572
rect 21726 16532 21732 16544
rect 21784 16532 21790 16584
rect 21910 16572 21916 16584
rect 21871 16544 21916 16572
rect 21910 16532 21916 16544
rect 21968 16532 21974 16584
rect 22020 16581 22048 16612
rect 23290 16600 23296 16652
rect 23348 16640 23354 16652
rect 24765 16643 24823 16649
rect 24765 16640 24777 16643
rect 23348 16612 24777 16640
rect 23348 16600 23354 16612
rect 24765 16609 24777 16612
rect 24811 16609 24823 16643
rect 28350 16640 28356 16652
rect 28311 16612 28356 16640
rect 24765 16603 24823 16609
rect 28350 16600 28356 16612
rect 28408 16600 28414 16652
rect 22005 16575 22063 16581
rect 22005 16541 22017 16575
rect 22051 16541 22063 16575
rect 22005 16535 22063 16541
rect 22097 16575 22155 16581
rect 22097 16541 22109 16575
rect 22143 16572 22155 16575
rect 22462 16572 22468 16584
rect 22143 16544 22468 16572
rect 22143 16541 22155 16544
rect 22097 16535 22155 16541
rect 22462 16532 22468 16544
rect 22520 16532 22526 16584
rect 23014 16532 23020 16584
rect 23072 16572 23078 16584
rect 23201 16575 23259 16581
rect 23201 16572 23213 16575
rect 23072 16544 23213 16572
rect 23072 16532 23078 16544
rect 23201 16541 23213 16544
rect 23247 16541 23259 16575
rect 23382 16572 23388 16584
rect 23343 16544 23388 16572
rect 23201 16535 23259 16541
rect 23382 16532 23388 16544
rect 23440 16532 23446 16584
rect 23477 16575 23535 16581
rect 23477 16541 23489 16575
rect 23523 16541 23535 16575
rect 23477 16535 23535 16541
rect 20714 16504 20720 16516
rect 20675 16476 20720 16504
rect 20714 16464 20720 16476
rect 20772 16464 20778 16516
rect 21174 16504 21180 16516
rect 21135 16476 21180 16504
rect 21174 16464 21180 16476
rect 21232 16464 21238 16516
rect 21361 16507 21419 16513
rect 21361 16473 21373 16507
rect 21407 16504 21419 16507
rect 22186 16504 22192 16516
rect 21407 16476 22192 16504
rect 21407 16473 21419 16476
rect 21361 16467 21419 16473
rect 22186 16464 22192 16476
rect 22244 16504 22250 16516
rect 22554 16504 22560 16516
rect 22244 16476 22560 16504
rect 22244 16464 22250 16476
rect 22554 16464 22560 16476
rect 22612 16464 22618 16516
rect 22833 16507 22891 16513
rect 22833 16473 22845 16507
rect 22879 16504 22891 16507
rect 23106 16504 23112 16516
rect 22879 16476 23112 16504
rect 22879 16473 22891 16476
rect 22833 16467 22891 16473
rect 23106 16464 23112 16476
rect 23164 16504 23170 16516
rect 23492 16504 23520 16535
rect 23566 16532 23572 16584
rect 23624 16572 23630 16584
rect 25038 16572 25044 16584
rect 23624 16544 25044 16572
rect 23624 16532 23630 16544
rect 25038 16532 25044 16544
rect 25096 16532 25102 16584
rect 23164 16476 23520 16504
rect 23164 16464 23170 16476
rect 23750 16464 23756 16516
rect 23808 16504 23814 16516
rect 24397 16507 24455 16513
rect 24397 16504 24409 16507
rect 23808 16476 24409 16504
rect 23808 16464 23814 16476
rect 24397 16473 24409 16476
rect 24443 16473 24455 16507
rect 24578 16504 24584 16516
rect 24539 16476 24584 16504
rect 24397 16467 24455 16473
rect 24578 16464 24584 16476
rect 24636 16464 24642 16516
rect 18892 16408 19656 16436
rect 19797 16439 19855 16445
rect 18785 16399 18843 16405
rect 19797 16405 19809 16439
rect 19843 16436 19855 16439
rect 19886 16436 19892 16448
rect 19843 16408 19892 16436
rect 19843 16405 19855 16408
rect 19797 16399 19855 16405
rect 19886 16396 19892 16408
rect 19944 16396 19950 16448
rect 20993 16439 21051 16445
rect 20993 16405 21005 16439
rect 21039 16436 21051 16439
rect 21082 16436 21088 16448
rect 21039 16408 21088 16436
rect 21039 16405 21051 16408
rect 20993 16399 21051 16405
rect 21082 16396 21088 16408
rect 21140 16396 21146 16448
rect 22373 16439 22431 16445
rect 22373 16405 22385 16439
rect 22419 16436 22431 16439
rect 23658 16436 23664 16448
rect 22419 16408 23664 16436
rect 22419 16405 22431 16408
rect 22373 16399 22431 16405
rect 23658 16396 23664 16408
rect 23716 16396 23722 16448
rect 1104 16346 28888 16368
rect 1104 16294 10214 16346
rect 10266 16294 10278 16346
rect 10330 16294 10342 16346
rect 10394 16294 10406 16346
rect 10458 16294 10470 16346
rect 10522 16294 19478 16346
rect 19530 16294 19542 16346
rect 19594 16294 19606 16346
rect 19658 16294 19670 16346
rect 19722 16294 19734 16346
rect 19786 16294 28888 16346
rect 1104 16272 28888 16294
rect 7650 16232 7656 16244
rect 7611 16204 7656 16232
rect 7650 16192 7656 16204
rect 7708 16192 7714 16244
rect 9306 16192 9312 16244
rect 9364 16232 9370 16244
rect 11882 16232 11888 16244
rect 9364 16204 11888 16232
rect 9364 16192 9370 16204
rect 11882 16192 11888 16204
rect 11940 16192 11946 16244
rect 11974 16192 11980 16244
rect 12032 16232 12038 16244
rect 12831 16235 12889 16241
rect 12831 16232 12843 16235
rect 12032 16204 12843 16232
rect 12032 16192 12038 16204
rect 12831 16201 12843 16204
rect 12877 16232 12889 16235
rect 12877 16204 13508 16232
rect 12877 16201 12889 16204
rect 12831 16195 12889 16201
rect 9766 16164 9772 16176
rect 8772 16136 9772 16164
rect 5813 16099 5871 16105
rect 5813 16065 5825 16099
rect 5859 16096 5871 16099
rect 5902 16096 5908 16108
rect 5859 16068 5908 16096
rect 5859 16065 5871 16068
rect 5813 16059 5871 16065
rect 5902 16056 5908 16068
rect 5960 16056 5966 16108
rect 5997 16099 6055 16105
rect 5997 16065 6009 16099
rect 6043 16096 6055 16099
rect 6638 16096 6644 16108
rect 6043 16068 6644 16096
rect 6043 16065 6055 16068
rect 5997 16059 6055 16065
rect 6638 16056 6644 16068
rect 6696 16056 6702 16108
rect 8772 16105 8800 16136
rect 9766 16124 9772 16136
rect 9824 16124 9830 16176
rect 12621 16167 12679 16173
rect 12621 16164 12633 16167
rect 11900 16136 12633 16164
rect 8757 16099 8815 16105
rect 6811 16089 6869 16095
rect 6811 16055 6823 16089
rect 6857 16055 6869 16089
rect 8757 16065 8769 16099
rect 8803 16065 8815 16099
rect 8757 16059 8815 16065
rect 8849 16099 8907 16105
rect 8849 16065 8861 16099
rect 8895 16096 8907 16099
rect 9214 16096 9220 16108
rect 8895 16068 9220 16096
rect 8895 16065 8907 16068
rect 8849 16059 8907 16065
rect 9214 16056 9220 16068
rect 9272 16056 9278 16108
rect 9582 16105 9588 16108
rect 9576 16059 9588 16105
rect 9640 16096 9646 16108
rect 11149 16099 11207 16105
rect 9640 16068 9676 16096
rect 9582 16056 9588 16059
rect 9640 16056 9646 16068
rect 11149 16065 11161 16099
rect 11195 16096 11207 16099
rect 11238 16096 11244 16108
rect 11195 16068 11244 16096
rect 11195 16065 11207 16068
rect 11149 16059 11207 16065
rect 11238 16056 11244 16068
rect 11296 16096 11302 16108
rect 11422 16096 11428 16108
rect 11296 16068 11428 16096
rect 11296 16056 11302 16068
rect 11422 16056 11428 16068
rect 11480 16056 11486 16108
rect 11698 16056 11704 16108
rect 11756 16096 11762 16108
rect 11900 16105 11928 16136
rect 12621 16133 12633 16136
rect 12667 16133 12679 16167
rect 13262 16164 13268 16176
rect 13223 16136 13268 16164
rect 12621 16127 12679 16133
rect 13262 16124 13268 16136
rect 13320 16124 13326 16176
rect 13480 16164 13508 16204
rect 13740 16204 14412 16232
rect 13538 16164 13544 16176
rect 13480 16133 13544 16164
rect 11885 16099 11943 16105
rect 13480 16102 13507 16133
rect 11885 16096 11897 16099
rect 11756 16068 11897 16096
rect 11756 16056 11762 16068
rect 11885 16065 11897 16068
rect 11931 16065 11943 16099
rect 13495 16099 13507 16102
rect 13541 16124 13544 16133
rect 13596 16124 13602 16176
rect 13541 16099 13553 16124
rect 13495 16093 13553 16099
rect 11885 16059 11943 16065
rect 6811 16049 6869 16055
rect 6831 15960 6859 16049
rect 7745 16031 7803 16037
rect 7745 15997 7757 16031
rect 7791 15997 7803 16031
rect 7745 15991 7803 15997
rect 7285 15963 7343 15969
rect 7285 15960 7297 15963
rect 6831 15932 7297 15960
rect 7285 15929 7297 15932
rect 7331 15929 7343 15963
rect 7285 15923 7343 15929
rect 7650 15920 7656 15972
rect 7708 15960 7714 15972
rect 7760 15960 7788 15991
rect 7834 15988 7840 16040
rect 7892 16028 7898 16040
rect 9306 16028 9312 16040
rect 7892 16000 7937 16028
rect 9267 16000 9312 16028
rect 7892 15988 7898 16000
rect 9306 15988 9312 16000
rect 9364 15988 9370 16040
rect 11977 16031 12035 16037
rect 11977 16028 11989 16031
rect 10336 16000 11989 16028
rect 7708 15932 9352 15960
rect 7708 15920 7714 15932
rect 5166 15852 5172 15904
rect 5224 15892 5230 15904
rect 5629 15895 5687 15901
rect 5629 15892 5641 15895
rect 5224 15864 5641 15892
rect 5224 15852 5230 15864
rect 5629 15861 5641 15864
rect 5675 15861 5687 15895
rect 5629 15855 5687 15861
rect 7009 15895 7067 15901
rect 7009 15861 7021 15895
rect 7055 15892 7067 15895
rect 8478 15892 8484 15904
rect 7055 15864 8484 15892
rect 7055 15861 7067 15864
rect 7009 15855 7067 15861
rect 8478 15852 8484 15864
rect 8536 15852 8542 15904
rect 9030 15892 9036 15904
rect 8991 15864 9036 15892
rect 9030 15852 9036 15864
rect 9088 15852 9094 15904
rect 9324 15892 9352 15932
rect 10336 15892 10364 16000
rect 11977 15997 11989 16000
rect 12023 15997 12035 16031
rect 11977 15991 12035 15997
rect 12069 16031 12127 16037
rect 12069 15997 12081 16031
rect 12115 16028 12127 16031
rect 12250 16028 12256 16040
rect 12115 16000 12256 16028
rect 12115 15997 12127 16000
rect 12069 15991 12127 15997
rect 11146 15920 11152 15972
rect 11204 15960 11210 15972
rect 12084 15960 12112 15991
rect 12250 15988 12256 16000
rect 12308 15988 12314 16040
rect 13740 16028 13768 16204
rect 13906 16124 13912 16176
rect 13964 16164 13970 16176
rect 13964 16136 14320 16164
rect 13964 16124 13970 16136
rect 13998 16096 14004 16108
rect 13959 16068 14004 16096
rect 13998 16056 14004 16068
rect 14056 16056 14062 16108
rect 14292 16105 14320 16136
rect 14384 16105 14412 16204
rect 15470 16192 15476 16244
rect 15528 16232 15534 16244
rect 16761 16235 16819 16241
rect 15528 16204 16528 16232
rect 15528 16192 15534 16204
rect 14458 16124 14464 16176
rect 14516 16164 14522 16176
rect 16500 16164 16528 16204
rect 16761 16201 16773 16235
rect 16807 16232 16819 16235
rect 16942 16232 16948 16244
rect 16807 16204 16948 16232
rect 16807 16201 16819 16204
rect 16761 16195 16819 16201
rect 16942 16192 16948 16204
rect 17000 16192 17006 16244
rect 17770 16232 17776 16244
rect 17236 16204 17776 16232
rect 16666 16164 16672 16176
rect 14516 16136 14872 16164
rect 16500 16136 16672 16164
rect 14516 16124 14522 16136
rect 14277 16099 14335 16105
rect 14277 16065 14289 16099
rect 14323 16065 14335 16099
rect 14277 16059 14335 16065
rect 14369 16099 14427 16105
rect 14369 16065 14381 16099
rect 14415 16065 14427 16099
rect 14550 16096 14556 16108
rect 14511 16068 14556 16096
rect 14369 16059 14427 16065
rect 14550 16056 14556 16068
rect 14608 16056 14614 16108
rect 14844 16105 14872 16136
rect 16666 16124 16672 16136
rect 16724 16164 16730 16176
rect 17037 16167 17095 16173
rect 17037 16164 17049 16167
rect 16724 16136 17049 16164
rect 16724 16124 16730 16136
rect 17037 16133 17049 16136
rect 17083 16133 17095 16167
rect 17037 16127 17095 16133
rect 14829 16099 14887 16105
rect 14829 16065 14841 16099
rect 14875 16065 14887 16099
rect 15102 16096 15108 16108
rect 15063 16068 15108 16096
rect 14829 16059 14887 16065
rect 15102 16056 15108 16068
rect 15160 16056 15166 16108
rect 15194 16056 15200 16108
rect 15252 16096 15258 16108
rect 16022 16096 16028 16108
rect 15252 16068 15297 16096
rect 15983 16068 16028 16096
rect 15252 16056 15258 16068
rect 16022 16056 16028 16068
rect 16080 16056 16086 16108
rect 16301 16099 16359 16105
rect 16301 16065 16313 16099
rect 16347 16096 16359 16099
rect 16482 16096 16488 16108
rect 16347 16068 16488 16096
rect 16347 16065 16359 16068
rect 16301 16059 16359 16065
rect 16482 16056 16488 16068
rect 16540 16056 16546 16108
rect 17236 16105 17264 16204
rect 17770 16192 17776 16204
rect 17828 16232 17834 16244
rect 19150 16232 19156 16244
rect 17828 16204 19156 16232
rect 17828 16192 17834 16204
rect 19150 16192 19156 16204
rect 19208 16192 19214 16244
rect 19334 16192 19340 16244
rect 19392 16232 19398 16244
rect 20257 16235 20315 16241
rect 20257 16232 20269 16235
rect 19392 16204 20269 16232
rect 19392 16192 19398 16204
rect 20257 16201 20269 16204
rect 20303 16201 20315 16235
rect 20257 16195 20315 16201
rect 21174 16192 21180 16244
rect 21232 16232 21238 16244
rect 24578 16232 24584 16244
rect 21232 16204 24584 16232
rect 21232 16192 21238 16204
rect 24578 16192 24584 16204
rect 24636 16232 24642 16244
rect 25317 16235 25375 16241
rect 25317 16232 25329 16235
rect 24636 16204 25329 16232
rect 24636 16192 24642 16204
rect 25317 16201 25329 16204
rect 25363 16201 25375 16235
rect 25317 16195 25375 16201
rect 17310 16124 17316 16176
rect 17368 16164 17374 16176
rect 19429 16167 19487 16173
rect 19429 16164 19441 16167
rect 17368 16136 19441 16164
rect 17368 16124 17374 16136
rect 17420 16105 17448 16136
rect 19429 16133 19441 16136
rect 19475 16164 19487 16167
rect 22462 16164 22468 16176
rect 19475 16136 20024 16164
rect 19475 16133 19487 16136
rect 19429 16127 19487 16133
rect 17221 16099 17279 16105
rect 17221 16065 17233 16099
rect 17267 16065 17279 16099
rect 17221 16059 17279 16065
rect 17405 16099 17463 16105
rect 17405 16065 17417 16099
rect 17451 16065 17463 16099
rect 17405 16059 17463 16065
rect 17589 16099 17647 16105
rect 17589 16065 17601 16099
rect 17635 16065 17647 16099
rect 17862 16096 17868 16108
rect 17823 16068 17868 16096
rect 17589 16059 17647 16065
rect 13004 16000 13768 16028
rect 14093 16031 14151 16037
rect 13004 15969 13032 16000
rect 14093 15997 14105 16031
rect 14139 16028 14151 16031
rect 14921 16031 14979 16037
rect 14921 16028 14933 16031
rect 14139 16000 14933 16028
rect 14139 15997 14151 16000
rect 14093 15991 14151 15997
rect 14921 15997 14933 16000
rect 14967 16028 14979 16031
rect 15746 16028 15752 16040
rect 14967 16000 15752 16028
rect 14967 15997 14979 16000
rect 14921 15991 14979 15997
rect 15746 15988 15752 16000
rect 15804 16028 15810 16040
rect 16114 16028 16120 16040
rect 15804 16000 15884 16028
rect 16075 16000 16120 16028
rect 15804 15988 15810 16000
rect 11204 15932 12112 15960
rect 12989 15963 13047 15969
rect 11204 15920 11210 15932
rect 12989 15929 13001 15963
rect 13035 15929 13047 15963
rect 12989 15923 13047 15929
rect 13633 15963 13691 15969
rect 13633 15929 13645 15963
rect 13679 15960 13691 15963
rect 15010 15960 15016 15972
rect 13679 15932 15016 15960
rect 13679 15929 13691 15932
rect 13633 15923 13691 15929
rect 15010 15920 15016 15932
rect 15068 15920 15074 15972
rect 15378 15960 15384 15972
rect 15339 15932 15384 15960
rect 15378 15920 15384 15932
rect 15436 15920 15442 15972
rect 15856 15969 15884 16000
rect 16114 15988 16120 16000
rect 16172 15988 16178 16040
rect 16850 15988 16856 16040
rect 16908 16028 16914 16040
rect 17604 16028 17632 16059
rect 17862 16056 17868 16068
rect 17920 16056 17926 16108
rect 18322 16096 18328 16108
rect 18283 16068 18328 16096
rect 18322 16056 18328 16068
rect 18380 16056 18386 16108
rect 18782 16056 18788 16108
rect 18840 16096 18846 16108
rect 18877 16099 18935 16105
rect 18877 16096 18889 16099
rect 18840 16068 18889 16096
rect 18840 16056 18846 16068
rect 18877 16065 18889 16068
rect 18923 16065 18935 16099
rect 18877 16059 18935 16065
rect 19150 16056 19156 16108
rect 19208 16096 19214 16108
rect 19797 16099 19855 16105
rect 19797 16096 19809 16099
rect 19208 16068 19809 16096
rect 19208 16056 19214 16068
rect 19797 16065 19809 16068
rect 19843 16065 19855 16099
rect 19797 16059 19855 16065
rect 19886 16056 19892 16108
rect 19944 16096 19950 16108
rect 19996 16105 20024 16136
rect 20916 16136 22468 16164
rect 19981 16099 20039 16105
rect 19981 16096 19993 16099
rect 19944 16068 19993 16096
rect 19944 16056 19950 16068
rect 19981 16065 19993 16068
rect 20027 16065 20039 16099
rect 19981 16059 20039 16065
rect 20070 16056 20076 16108
rect 20128 16096 20134 16108
rect 20916 16105 20944 16136
rect 20901 16099 20959 16105
rect 20128 16068 20173 16096
rect 20128 16056 20134 16068
rect 20901 16065 20913 16099
rect 20947 16065 20959 16099
rect 20901 16059 20959 16065
rect 20993 16099 21051 16105
rect 20993 16065 21005 16099
rect 21039 16065 21051 16099
rect 20993 16059 21051 16065
rect 18969 16031 19027 16037
rect 16908 16000 18828 16028
rect 16908 15988 16914 16000
rect 15841 15963 15899 15969
rect 15841 15929 15853 15963
rect 15887 15929 15899 15963
rect 15841 15923 15899 15929
rect 15948 15932 18736 15960
rect 10686 15892 10692 15904
rect 9324 15864 10364 15892
rect 10647 15864 10692 15892
rect 10686 15852 10692 15864
rect 10744 15852 10750 15904
rect 10870 15852 10876 15904
rect 10928 15892 10934 15904
rect 10965 15895 11023 15901
rect 10965 15892 10977 15895
rect 10928 15864 10977 15892
rect 10928 15852 10934 15864
rect 10965 15861 10977 15864
rect 11011 15861 11023 15895
rect 10965 15855 11023 15861
rect 11238 15852 11244 15904
rect 11296 15892 11302 15904
rect 11517 15895 11575 15901
rect 11517 15892 11529 15895
rect 11296 15864 11529 15892
rect 11296 15852 11302 15864
rect 11517 15861 11529 15864
rect 11563 15861 11575 15895
rect 12802 15892 12808 15904
rect 12715 15864 12808 15892
rect 11517 15855 11575 15861
rect 12802 15852 12808 15864
rect 12860 15892 12866 15904
rect 13449 15895 13507 15901
rect 13449 15892 13461 15895
rect 12860 15864 13461 15892
rect 12860 15852 12866 15864
rect 13449 15861 13461 15864
rect 13495 15892 13507 15895
rect 13538 15892 13544 15904
rect 13495 15864 13544 15892
rect 13495 15861 13507 15864
rect 13449 15855 13507 15861
rect 13538 15852 13544 15864
rect 13596 15892 13602 15904
rect 15948 15892 15976 15932
rect 13596 15864 15976 15892
rect 16301 15895 16359 15901
rect 13596 15852 13602 15864
rect 16301 15861 16313 15895
rect 16347 15892 16359 15895
rect 17770 15892 17776 15904
rect 16347 15864 17776 15892
rect 16347 15861 16359 15864
rect 16301 15855 16359 15861
rect 17770 15852 17776 15864
rect 17828 15852 17834 15904
rect 18708 15901 18736 15932
rect 18693 15895 18751 15901
rect 18693 15861 18705 15895
rect 18739 15861 18751 15895
rect 18800 15892 18828 16000
rect 18969 15997 18981 16031
rect 19015 16028 19027 16031
rect 20346 16028 20352 16040
rect 19015 16000 20352 16028
rect 19015 15997 19027 16000
rect 18969 15991 19027 15997
rect 20346 15988 20352 16000
rect 20404 15988 20410 16040
rect 21008 15972 21036 16059
rect 21082 16056 21088 16108
rect 21140 16096 21146 16108
rect 21269 16099 21327 16105
rect 21140 16068 21185 16096
rect 21140 16056 21146 16068
rect 21269 16065 21281 16099
rect 21315 16096 21327 16099
rect 21726 16096 21732 16108
rect 21315 16068 21732 16096
rect 21315 16065 21327 16068
rect 21269 16059 21327 16065
rect 21284 16028 21312 16059
rect 21726 16056 21732 16068
rect 21784 16096 21790 16108
rect 21821 16099 21879 16105
rect 21821 16096 21833 16099
rect 21784 16068 21833 16096
rect 21784 16056 21790 16068
rect 21821 16065 21833 16068
rect 21867 16065 21879 16099
rect 22002 16096 22008 16108
rect 21963 16068 22008 16096
rect 21821 16059 21879 16065
rect 22002 16056 22008 16068
rect 22060 16056 22066 16108
rect 22097 16099 22155 16105
rect 22097 16065 22109 16099
rect 22143 16065 22155 16099
rect 22097 16059 22155 16065
rect 22189 16099 22247 16105
rect 22189 16065 22201 16099
rect 22235 16096 22247 16099
rect 22296 16096 22324 16136
rect 22462 16124 22468 16136
rect 22520 16124 22526 16176
rect 23661 16167 23719 16173
rect 23661 16133 23673 16167
rect 23707 16164 23719 16167
rect 24182 16167 24240 16173
rect 24182 16164 24194 16167
rect 23707 16136 24194 16164
rect 23707 16133 23719 16136
rect 23661 16127 23719 16133
rect 24182 16133 24194 16136
rect 24228 16133 24240 16167
rect 24182 16127 24240 16133
rect 23014 16096 23020 16108
rect 22235 16068 22324 16096
rect 22975 16068 23020 16096
rect 22235 16065 22247 16068
rect 22189 16059 22247 16065
rect 21100 16000 21312 16028
rect 21100 15972 21128 16000
rect 22112 15972 22140 16059
rect 23014 16056 23020 16068
rect 23072 16056 23078 16108
rect 23198 16105 23204 16108
rect 23196 16096 23204 16105
rect 23159 16068 23204 16096
rect 23196 16059 23204 16068
rect 23198 16056 23204 16059
rect 23256 16056 23262 16108
rect 23296 16099 23354 16105
rect 23296 16065 23308 16099
rect 23342 16065 23354 16099
rect 23296 16059 23354 16065
rect 19426 15960 19432 15972
rect 19387 15932 19432 15960
rect 19426 15920 19432 15932
rect 19484 15920 19490 15972
rect 20990 15920 20996 15972
rect 21048 15920 21054 15972
rect 21082 15920 21088 15972
rect 21140 15920 21146 15972
rect 22094 15920 22100 15972
rect 22152 15920 22158 15972
rect 23106 15920 23112 15972
rect 23164 15960 23170 15972
rect 23311 15960 23339 16059
rect 23382 16056 23388 16108
rect 23440 16096 23446 16108
rect 25593 16099 25651 16105
rect 25593 16096 25605 16099
rect 23440 16068 25605 16096
rect 23440 16056 23446 16068
rect 25593 16065 25605 16068
rect 25639 16096 25651 16099
rect 26418 16096 26424 16108
rect 25639 16068 26424 16096
rect 25639 16065 25651 16068
rect 25593 16059 25651 16065
rect 26418 16056 26424 16068
rect 26476 16056 26482 16108
rect 23934 16028 23940 16040
rect 23895 16000 23940 16028
rect 23934 15988 23940 16000
rect 23992 15988 23998 16040
rect 23164 15932 23339 15960
rect 23164 15920 23170 15932
rect 19797 15895 19855 15901
rect 19797 15892 19809 15895
rect 18800 15864 19809 15892
rect 18693 15855 18751 15861
rect 19797 15861 19809 15864
rect 19843 15892 19855 15895
rect 19886 15892 19892 15904
rect 19843 15864 19892 15892
rect 19843 15861 19855 15864
rect 19797 15855 19855 15861
rect 19886 15852 19892 15864
rect 19944 15852 19950 15904
rect 20625 15895 20683 15901
rect 20625 15861 20637 15895
rect 20671 15892 20683 15895
rect 21542 15892 21548 15904
rect 20671 15864 21548 15892
rect 20671 15861 20683 15864
rect 20625 15855 20683 15861
rect 21542 15852 21548 15864
rect 21600 15852 21606 15904
rect 22465 15895 22523 15901
rect 22465 15861 22477 15895
rect 22511 15892 22523 15895
rect 22830 15892 22836 15904
rect 22511 15864 22836 15892
rect 22511 15861 22523 15864
rect 22465 15855 22523 15861
rect 22830 15852 22836 15864
rect 22888 15852 22894 15904
rect 1104 15802 28888 15824
rect 1104 15750 5582 15802
rect 5634 15750 5646 15802
rect 5698 15750 5710 15802
rect 5762 15750 5774 15802
rect 5826 15750 5838 15802
rect 5890 15750 14846 15802
rect 14898 15750 14910 15802
rect 14962 15750 14974 15802
rect 15026 15750 15038 15802
rect 15090 15750 15102 15802
rect 15154 15750 24110 15802
rect 24162 15750 24174 15802
rect 24226 15750 24238 15802
rect 24290 15750 24302 15802
rect 24354 15750 24366 15802
rect 24418 15750 28888 15802
rect 1104 15728 28888 15750
rect 5902 15648 5908 15700
rect 5960 15688 5966 15700
rect 7285 15691 7343 15697
rect 7285 15688 7297 15691
rect 5960 15660 7297 15688
rect 5960 15648 5966 15660
rect 7285 15657 7297 15660
rect 7331 15657 7343 15691
rect 8294 15688 8300 15700
rect 8255 15660 8300 15688
rect 7285 15651 7343 15657
rect 8294 15648 8300 15660
rect 8352 15648 8358 15700
rect 9582 15648 9588 15700
rect 9640 15688 9646 15700
rect 9677 15691 9735 15697
rect 9677 15688 9689 15691
rect 9640 15660 9689 15688
rect 9640 15648 9646 15660
rect 9677 15657 9689 15660
rect 9723 15657 9735 15691
rect 11698 15688 11704 15700
rect 11659 15660 11704 15688
rect 9677 15651 9735 15657
rect 11698 15648 11704 15660
rect 11756 15648 11762 15700
rect 11882 15648 11888 15700
rect 11940 15688 11946 15700
rect 13538 15688 13544 15700
rect 11940 15660 13124 15688
rect 13499 15660 13544 15688
rect 11940 15648 11946 15660
rect 7009 15623 7067 15629
rect 7009 15589 7021 15623
rect 7055 15620 7067 15623
rect 7650 15620 7656 15632
rect 7055 15592 7656 15620
rect 7055 15589 7067 15592
rect 7009 15583 7067 15589
rect 7650 15580 7656 15592
rect 7708 15580 7714 15632
rect 7282 15512 7288 15564
rect 7340 15552 7346 15564
rect 7834 15552 7840 15564
rect 7340 15524 7840 15552
rect 7340 15512 7346 15524
rect 7834 15512 7840 15524
rect 7892 15512 7898 15564
rect 10870 15512 10876 15564
rect 10928 15552 10934 15564
rect 13096 15561 13124 15660
rect 13538 15648 13544 15660
rect 13596 15648 13602 15700
rect 13725 15691 13783 15697
rect 13725 15657 13737 15691
rect 13771 15688 13783 15691
rect 15194 15688 15200 15700
rect 13771 15660 15200 15688
rect 13771 15657 13783 15660
rect 13725 15651 13783 15657
rect 15194 15648 15200 15660
rect 15252 15648 15258 15700
rect 22002 15648 22008 15700
rect 22060 15688 22066 15700
rect 22097 15691 22155 15697
rect 22097 15688 22109 15691
rect 22060 15660 22109 15688
rect 22060 15648 22066 15660
rect 22097 15657 22109 15660
rect 22143 15657 22155 15691
rect 22097 15651 22155 15657
rect 22186 15648 22192 15700
rect 22244 15688 22250 15700
rect 22922 15688 22928 15700
rect 22244 15660 22928 15688
rect 22244 15648 22250 15660
rect 22922 15648 22928 15660
rect 22980 15688 22986 15700
rect 22980 15660 23520 15688
rect 22980 15648 22986 15660
rect 20530 15620 20536 15632
rect 20491 15592 20536 15620
rect 20530 15580 20536 15592
rect 20588 15580 20594 15632
rect 21085 15623 21143 15629
rect 21085 15589 21097 15623
rect 21131 15620 21143 15623
rect 22462 15620 22468 15632
rect 21131 15592 22468 15620
rect 21131 15589 21143 15592
rect 21085 15583 21143 15589
rect 22462 15580 22468 15592
rect 22520 15580 22526 15632
rect 23014 15580 23020 15632
rect 23072 15580 23078 15632
rect 23198 15580 23204 15632
rect 23256 15620 23262 15632
rect 23256 15592 23336 15620
rect 23256 15580 23262 15592
rect 11057 15555 11115 15561
rect 11057 15552 11069 15555
rect 10928 15524 11069 15552
rect 10928 15512 10934 15524
rect 11057 15521 11069 15524
rect 11103 15521 11115 15555
rect 11057 15515 11115 15521
rect 13081 15555 13139 15561
rect 13081 15521 13093 15555
rect 13127 15552 13139 15555
rect 14093 15555 14151 15561
rect 14093 15552 14105 15555
rect 13127 15524 14105 15552
rect 13127 15521 13139 15524
rect 13081 15515 13139 15521
rect 14093 15521 14105 15524
rect 14139 15521 14151 15555
rect 17862 15552 17868 15564
rect 17823 15524 17868 15552
rect 14093 15515 14151 15521
rect 17862 15512 17868 15524
rect 17920 15552 17926 15564
rect 19426 15552 19432 15564
rect 17920 15524 19432 15552
rect 17920 15512 17926 15524
rect 19426 15512 19432 15524
rect 19484 15552 19490 15564
rect 19521 15555 19579 15561
rect 19521 15552 19533 15555
rect 19484 15524 19533 15552
rect 19484 15512 19490 15524
rect 19521 15521 19533 15524
rect 19567 15521 19579 15555
rect 20346 15552 20352 15564
rect 20259 15524 20352 15552
rect 19521 15515 19579 15521
rect 20346 15512 20352 15524
rect 20404 15552 20410 15564
rect 21450 15552 21456 15564
rect 20404 15524 21456 15552
rect 20404 15512 20410 15524
rect 21450 15512 21456 15524
rect 21508 15512 21514 15564
rect 23032 15552 23060 15580
rect 21836 15524 22600 15552
rect 23032 15524 23152 15552
rect 5166 15484 5172 15496
rect 5127 15456 5172 15484
rect 5166 15444 5172 15456
rect 5224 15444 5230 15496
rect 5626 15484 5632 15496
rect 5587 15456 5632 15484
rect 5626 15444 5632 15456
rect 5684 15444 5690 15496
rect 7650 15484 7656 15496
rect 7611 15456 7656 15484
rect 7650 15444 7656 15456
rect 7708 15444 7714 15496
rect 7742 15444 7748 15496
rect 7800 15484 7806 15496
rect 8478 15484 8484 15496
rect 7800 15456 7845 15484
rect 8439 15456 8484 15484
rect 7800 15444 7806 15456
rect 8478 15444 8484 15456
rect 8536 15444 8542 15496
rect 9030 15444 9036 15496
rect 9088 15484 9094 15496
rect 9493 15487 9551 15493
rect 9493 15484 9505 15487
rect 9088 15456 9505 15484
rect 9088 15444 9094 15456
rect 9493 15453 9505 15456
rect 9539 15453 9551 15487
rect 11238 15484 11244 15496
rect 11199 15456 11244 15484
rect 9493 15447 9551 15453
rect 11238 15444 11244 15456
rect 11296 15444 11302 15496
rect 15838 15484 15844 15496
rect 13587 15453 13645 15459
rect 15799 15456 15844 15484
rect 13587 15450 13599 15453
rect 5874 15419 5932 15425
rect 5874 15416 5886 15419
rect 5368 15388 5886 15416
rect 5368 15357 5396 15388
rect 5874 15385 5886 15388
rect 5920 15385 5932 15419
rect 5874 15379 5932 15385
rect 7190 15376 7196 15428
rect 7248 15416 7254 15428
rect 7760 15416 7788 15444
rect 7248 15388 7788 15416
rect 11425 15419 11483 15425
rect 7248 15376 7254 15388
rect 11425 15385 11437 15419
rect 11471 15416 11483 15419
rect 12342 15416 12348 15428
rect 11471 15388 12348 15416
rect 11471 15385 11483 15388
rect 11425 15379 11483 15385
rect 12342 15376 12348 15388
rect 12400 15376 12406 15428
rect 12526 15376 12532 15428
rect 12584 15416 12590 15428
rect 12814 15419 12872 15425
rect 12814 15416 12826 15419
rect 12584 15388 12826 15416
rect 12584 15376 12590 15388
rect 12814 15385 12826 15388
rect 12860 15385 12872 15419
rect 12814 15379 12872 15385
rect 13357 15419 13415 15425
rect 13357 15385 13369 15419
rect 13403 15385 13415 15419
rect 13572 15419 13599 15450
rect 13633 15428 13645 15453
rect 15838 15444 15844 15456
rect 15896 15444 15902 15496
rect 16022 15444 16028 15496
rect 16080 15484 16086 15496
rect 18141 15487 18199 15493
rect 18141 15484 18153 15487
rect 16080 15456 18153 15484
rect 16080 15444 16086 15456
rect 18141 15453 18153 15456
rect 18187 15453 18199 15487
rect 18141 15447 18199 15453
rect 18414 15444 18420 15496
rect 18472 15484 18478 15496
rect 19245 15487 19303 15493
rect 19245 15484 19257 15487
rect 18472 15456 19257 15484
rect 18472 15444 18478 15456
rect 19245 15453 19257 15456
rect 19291 15484 19303 15487
rect 20070 15484 20076 15496
rect 19291 15456 20076 15484
rect 19291 15453 19303 15456
rect 19245 15447 19303 15453
rect 20070 15444 20076 15456
rect 20128 15444 20134 15496
rect 21082 15444 21088 15496
rect 21140 15484 21146 15496
rect 21269 15487 21327 15493
rect 21269 15484 21281 15487
rect 21140 15456 21281 15484
rect 21140 15444 21146 15456
rect 21269 15453 21281 15456
rect 21315 15484 21327 15487
rect 21836 15484 21864 15524
rect 21315 15456 21864 15484
rect 21315 15453 21327 15456
rect 21269 15447 21327 15453
rect 22370 15444 22376 15496
rect 22428 15484 22434 15496
rect 22572 15493 22600 15524
rect 22557 15487 22615 15493
rect 22428 15456 22473 15484
rect 22428 15444 22434 15456
rect 22557 15453 22569 15487
rect 22603 15484 22615 15487
rect 22646 15484 22652 15496
rect 22603 15456 22652 15484
rect 22603 15453 22615 15456
rect 22557 15447 22615 15453
rect 22646 15444 22652 15456
rect 22704 15444 22710 15496
rect 23023 15487 23081 15493
rect 23023 15453 23035 15487
rect 23069 15486 23081 15487
rect 23124 15486 23152 15524
rect 23308 15493 23336 15592
rect 23293 15487 23351 15493
rect 23069 15458 23152 15486
rect 23196 15481 23254 15487
rect 23069 15453 23081 15458
rect 23023 15447 23081 15453
rect 23196 15447 23208 15481
rect 23242 15447 23254 15481
rect 23293 15453 23305 15487
rect 23339 15453 23351 15487
rect 23293 15447 23351 15453
rect 23405 15487 23463 15493
rect 23405 15453 23417 15487
rect 23451 15484 23463 15487
rect 23492 15484 23520 15660
rect 23842 15648 23848 15700
rect 23900 15688 23906 15700
rect 24029 15691 24087 15697
rect 24029 15688 24041 15691
rect 23900 15660 24041 15688
rect 23900 15648 23906 15660
rect 24029 15657 24041 15660
rect 24075 15688 24087 15691
rect 28166 15688 28172 15700
rect 24075 15660 28172 15688
rect 24075 15657 24087 15660
rect 24029 15651 24087 15657
rect 28166 15648 28172 15660
rect 28224 15648 28230 15700
rect 23934 15512 23940 15564
rect 23992 15552 23998 15564
rect 24397 15555 24455 15561
rect 24397 15552 24409 15555
rect 23992 15524 24409 15552
rect 23992 15512 23998 15524
rect 24397 15521 24409 15524
rect 24443 15521 24455 15555
rect 24397 15515 24455 15521
rect 25130 15484 25136 15496
rect 23451 15456 25136 15484
rect 23451 15453 23463 15456
rect 23405 15447 23463 15453
rect 23196 15441 23254 15447
rect 25130 15444 25136 15456
rect 25188 15444 25194 15496
rect 28350 15484 28356 15496
rect 28311 15456 28356 15484
rect 28350 15444 28356 15456
rect 28408 15444 28414 15496
rect 13633 15419 13636 15428
rect 13572 15388 13636 15419
rect 13357 15379 13415 15385
rect 5353 15351 5411 15357
rect 5353 15317 5365 15351
rect 5399 15317 5411 15351
rect 5353 15311 5411 15317
rect 10686 15308 10692 15360
rect 10744 15348 10750 15360
rect 13372 15348 13400 15379
rect 13630 15376 13636 15388
rect 13688 15376 13694 15428
rect 14360 15419 14418 15425
rect 14360 15385 14372 15419
rect 14406 15416 14418 15419
rect 15010 15416 15016 15428
rect 14406 15388 15016 15416
rect 14406 15385 14418 15388
rect 14360 15379 14418 15385
rect 15010 15376 15016 15388
rect 15068 15376 15074 15428
rect 20714 15376 20720 15428
rect 20772 15416 20778 15428
rect 20809 15419 20867 15425
rect 20809 15416 20821 15419
rect 20772 15388 20821 15416
rect 20772 15376 20778 15388
rect 20809 15385 20821 15388
rect 20855 15385 20867 15419
rect 20809 15379 20867 15385
rect 21729 15419 21787 15425
rect 21729 15385 21741 15419
rect 21775 15385 21787 15419
rect 21910 15416 21916 15428
rect 21871 15388 21916 15416
rect 21729 15379 21787 15385
rect 10744 15320 13400 15348
rect 10744 15308 10750 15320
rect 14090 15308 14096 15360
rect 14148 15348 14154 15360
rect 14642 15348 14648 15360
rect 14148 15320 14648 15348
rect 14148 15308 14154 15320
rect 14642 15308 14648 15320
rect 14700 15308 14706 15360
rect 15378 15308 15384 15360
rect 15436 15348 15442 15360
rect 15473 15351 15531 15357
rect 15473 15348 15485 15351
rect 15436 15320 15485 15348
rect 15436 15308 15442 15320
rect 15473 15317 15485 15320
rect 15519 15317 15531 15351
rect 17126 15348 17132 15360
rect 17087 15320 17132 15348
rect 15473 15311 15531 15317
rect 17126 15308 17132 15320
rect 17184 15308 17190 15360
rect 21744 15348 21772 15379
rect 21910 15376 21916 15388
rect 21968 15376 21974 15428
rect 22554 15348 22560 15360
rect 21744 15320 22560 15348
rect 22554 15308 22560 15320
rect 22612 15308 22618 15360
rect 22741 15351 22799 15357
rect 22741 15317 22753 15351
rect 22787 15348 22799 15351
rect 22922 15348 22928 15360
rect 22787 15320 22928 15348
rect 22787 15317 22799 15320
rect 22741 15311 22799 15317
rect 22922 15308 22928 15320
rect 22980 15308 22986 15360
rect 23216 15348 23244 15441
rect 23566 15416 23572 15428
rect 23400 15388 23572 15416
rect 23400 15348 23428 15388
rect 23566 15376 23572 15388
rect 23624 15376 23630 15428
rect 23661 15419 23719 15425
rect 23661 15385 23673 15419
rect 23707 15416 23719 15419
rect 24642 15419 24700 15425
rect 24642 15416 24654 15419
rect 23707 15388 24654 15416
rect 23707 15385 23719 15388
rect 23661 15379 23719 15385
rect 24642 15385 24654 15388
rect 24688 15385 24700 15419
rect 24642 15379 24700 15385
rect 23216 15320 23428 15348
rect 23934 15308 23940 15360
rect 23992 15348 23998 15360
rect 25777 15351 25835 15357
rect 25777 15348 25789 15351
rect 23992 15320 25789 15348
rect 23992 15308 23998 15320
rect 25777 15317 25789 15320
rect 25823 15317 25835 15351
rect 25777 15311 25835 15317
rect 1104 15258 28888 15280
rect 1104 15206 10214 15258
rect 10266 15206 10278 15258
rect 10330 15206 10342 15258
rect 10394 15206 10406 15258
rect 10458 15206 10470 15258
rect 10522 15206 19478 15258
rect 19530 15206 19542 15258
rect 19594 15206 19606 15258
rect 19658 15206 19670 15258
rect 19722 15206 19734 15258
rect 19786 15206 28888 15258
rect 1104 15184 28888 15206
rect 10873 15147 10931 15153
rect 10873 15113 10885 15147
rect 10919 15144 10931 15147
rect 11146 15144 11152 15156
rect 10919 15116 11152 15144
rect 10919 15113 10931 15116
rect 10873 15107 10931 15113
rect 11146 15104 11152 15116
rect 11204 15104 11210 15156
rect 12526 15144 12532 15156
rect 12487 15116 12532 15144
rect 12526 15104 12532 15116
rect 12584 15104 12590 15156
rect 15010 15144 15016 15156
rect 14971 15116 15016 15144
rect 15010 15104 15016 15116
rect 15068 15104 15074 15156
rect 16206 15144 16212 15156
rect 15672 15116 16212 15144
rect 8202 15036 8208 15088
rect 8260 15076 8266 15088
rect 9738 15079 9796 15085
rect 9738 15076 9750 15079
rect 8260 15048 9750 15076
rect 8260 15036 8266 15048
rect 9738 15045 9750 15048
rect 9784 15045 9796 15079
rect 9738 15039 9796 15045
rect 10594 15036 10600 15088
rect 10652 15076 10658 15088
rect 12805 15079 12863 15085
rect 12805 15076 12817 15079
rect 10652 15048 12817 15076
rect 10652 15036 10658 15048
rect 12805 15045 12817 15048
rect 12851 15076 12863 15079
rect 15562 15076 15568 15088
rect 12851 15048 15568 15076
rect 12851 15045 12863 15048
rect 12805 15039 12863 15045
rect 15562 15036 15568 15048
rect 15620 15036 15626 15088
rect 5626 14968 5632 15020
rect 5684 15008 5690 15020
rect 5994 15008 6000 15020
rect 5684 14980 6000 15008
rect 5684 14968 5690 14980
rect 5994 14968 6000 14980
rect 6052 15008 6058 15020
rect 8110 15017 8116 15020
rect 7837 15011 7895 15017
rect 7837 15008 7849 15011
rect 6052 14980 7849 15008
rect 6052 14968 6058 14980
rect 7837 14977 7849 14980
rect 7883 14977 7895 15011
rect 7837 14971 7895 14977
rect 8104 14971 8116 15017
rect 8168 15008 8174 15020
rect 8168 14980 8204 15008
rect 8110 14968 8116 14971
rect 8168 14968 8174 14980
rect 9306 14968 9312 15020
rect 9364 15008 9370 15020
rect 9493 15011 9551 15017
rect 9493 15008 9505 15011
rect 9364 14980 9505 15008
rect 9364 14968 9370 14980
rect 9493 14977 9505 14980
rect 9539 14977 9551 15011
rect 9493 14971 9551 14977
rect 11422 14968 11428 15020
rect 11480 15008 11486 15020
rect 11793 15011 11851 15017
rect 11793 15008 11805 15011
rect 11480 14980 11805 15008
rect 11480 14968 11486 14980
rect 11793 14977 11805 14980
rect 11839 15008 11851 15011
rect 11974 15008 11980 15020
rect 11839 14980 11980 15008
rect 11839 14977 11851 14980
rect 11793 14971 11851 14977
rect 11974 14968 11980 14980
rect 12032 14968 12038 15020
rect 12342 15008 12348 15020
rect 12303 14980 12348 15008
rect 12342 14968 12348 14980
rect 12400 14968 12406 15020
rect 13538 15008 13544 15020
rect 13499 14980 13544 15008
rect 13538 14968 13544 14980
rect 13596 14968 13602 15020
rect 13725 15011 13783 15017
rect 13725 14977 13737 15011
rect 13771 14977 13783 15011
rect 13725 14971 13783 14977
rect 13630 14900 13636 14952
rect 13688 14940 13694 14952
rect 13740 14940 13768 14971
rect 13906 14968 13912 15020
rect 13964 15008 13970 15020
rect 14274 15008 14280 15020
rect 13964 14980 14280 15008
rect 13964 14968 13970 14980
rect 14274 14968 14280 14980
rect 14332 14968 14338 15020
rect 15194 14968 15200 15020
rect 15252 15006 15258 15020
rect 15289 15011 15347 15017
rect 15289 15006 15301 15011
rect 15252 14978 15301 15006
rect 15252 14968 15258 14978
rect 15289 14977 15301 14978
rect 15335 14977 15347 15011
rect 15289 14971 15347 14977
rect 15381 15011 15439 15017
rect 15381 14977 15393 15011
rect 15427 14977 15439 15011
rect 15381 14971 15439 14977
rect 15396 14940 15424 14971
rect 15470 14968 15476 15020
rect 15528 15008 15534 15020
rect 15672 15017 15700 15116
rect 16206 15104 16212 15116
rect 16264 15104 16270 15156
rect 16301 15147 16359 15153
rect 16301 15113 16313 15147
rect 16347 15144 16359 15147
rect 16758 15144 16764 15156
rect 16347 15116 16764 15144
rect 16347 15113 16359 15116
rect 16301 15107 16359 15113
rect 16758 15104 16764 15116
rect 16816 15104 16822 15156
rect 17770 15144 17776 15156
rect 17731 15116 17776 15144
rect 17770 15104 17776 15116
rect 17828 15104 17834 15156
rect 19429 15147 19487 15153
rect 19429 15113 19441 15147
rect 19475 15144 19487 15147
rect 19889 15147 19947 15153
rect 19889 15144 19901 15147
rect 19475 15116 19901 15144
rect 19475 15113 19487 15116
rect 19429 15107 19487 15113
rect 19889 15113 19901 15116
rect 19935 15113 19947 15147
rect 20438 15144 20444 15156
rect 19889 15107 19947 15113
rect 20180 15116 20444 15144
rect 16022 15036 16028 15088
rect 16080 15076 16086 15088
rect 17788 15076 17816 15104
rect 16080 15048 17080 15076
rect 16080 15036 16086 15048
rect 15657 15011 15715 15017
rect 15528 14980 15573 15008
rect 15528 14968 15534 14980
rect 15657 14977 15669 15011
rect 15703 14977 15715 15011
rect 15657 14971 15715 14977
rect 16117 15011 16175 15017
rect 16117 14977 16129 15011
rect 16163 15008 16175 15011
rect 16206 15008 16212 15020
rect 16163 14980 16212 15008
rect 16163 14977 16175 14980
rect 16117 14971 16175 14977
rect 15746 14940 15752 14952
rect 13688 14912 15752 14940
rect 13688 14900 13694 14912
rect 15746 14900 15752 14912
rect 15804 14900 15810 14952
rect 12894 14832 12900 14884
rect 12952 14872 12958 14884
rect 14369 14875 14427 14881
rect 12952 14844 14320 14872
rect 12952 14832 12958 14844
rect 9217 14807 9275 14813
rect 9217 14773 9229 14807
rect 9263 14804 9275 14807
rect 9398 14804 9404 14816
rect 9263 14776 9404 14804
rect 9263 14773 9275 14776
rect 9217 14767 9275 14773
rect 9398 14764 9404 14776
rect 9456 14764 9462 14816
rect 11330 14764 11336 14816
rect 11388 14804 11394 14816
rect 11885 14807 11943 14813
rect 11885 14804 11897 14807
rect 11388 14776 11897 14804
rect 11388 14764 11394 14776
rect 11885 14773 11897 14776
rect 11931 14773 11943 14807
rect 13262 14804 13268 14816
rect 13223 14776 13268 14804
rect 11885 14767 11943 14773
rect 13262 14764 13268 14776
rect 13320 14764 13326 14816
rect 13633 14807 13691 14813
rect 13633 14773 13645 14807
rect 13679 14804 13691 14807
rect 14182 14804 14188 14816
rect 13679 14776 14188 14804
rect 13679 14773 13691 14776
rect 13633 14767 13691 14773
rect 14182 14764 14188 14776
rect 14240 14764 14246 14816
rect 14292 14804 14320 14844
rect 14369 14841 14381 14875
rect 14415 14872 14427 14875
rect 14458 14872 14464 14884
rect 14415 14844 14464 14872
rect 14415 14841 14427 14844
rect 14369 14835 14427 14841
rect 14458 14832 14464 14844
rect 14516 14832 14522 14884
rect 15838 14872 15844 14884
rect 14660 14844 15844 14872
rect 14660 14804 14688 14844
rect 15838 14832 15844 14844
rect 15896 14832 15902 14884
rect 16132 14872 16160 14971
rect 16206 14968 16212 14980
rect 16264 14968 16270 15020
rect 16301 15011 16359 15017
rect 16301 14977 16313 15011
rect 16347 14977 16359 15011
rect 16301 14971 16359 14977
rect 16040 14844 16160 14872
rect 16316 14872 16344 14971
rect 16482 14968 16488 15020
rect 16540 15008 16546 15020
rect 16761 15011 16819 15017
rect 16761 15008 16773 15011
rect 16540 14980 16773 15008
rect 16540 14968 16546 14980
rect 16761 14977 16773 14980
rect 16807 14977 16819 15011
rect 16761 14971 16819 14977
rect 16850 14968 16856 15020
rect 16908 15008 16914 15020
rect 16945 15011 17003 15017
rect 16945 15008 16957 15011
rect 16908 14980 16957 15008
rect 16908 14968 16914 14980
rect 16945 14977 16957 14980
rect 16991 14977 17003 15011
rect 16945 14971 17003 14977
rect 16390 14900 16396 14952
rect 16448 14940 16454 14952
rect 16669 14943 16727 14949
rect 16669 14940 16681 14943
rect 16448 14912 16681 14940
rect 16448 14900 16454 14912
rect 16669 14909 16681 14912
rect 16715 14909 16727 14943
rect 17052 14940 17080 15048
rect 17236 15048 17816 15076
rect 17236 15017 17264 15048
rect 19794 15036 19800 15088
rect 19852 15076 19858 15088
rect 20041 15079 20099 15085
rect 20041 15076 20053 15079
rect 19852 15048 20053 15076
rect 19852 15036 19858 15048
rect 20041 15045 20053 15048
rect 20087 15076 20099 15079
rect 20180 15076 20208 15116
rect 20438 15104 20444 15116
rect 20496 15104 20502 15156
rect 21266 15144 21272 15156
rect 21227 15116 21272 15144
rect 21266 15104 21272 15116
rect 21324 15104 21330 15156
rect 22002 15144 22008 15156
rect 21963 15116 22008 15144
rect 22002 15104 22008 15116
rect 22060 15104 22066 15156
rect 25130 15144 25136 15156
rect 25091 15116 25136 15144
rect 25130 15104 25136 15116
rect 25188 15104 25194 15156
rect 20087 15048 20208 15076
rect 20257 15079 20315 15085
rect 20087 15045 20099 15048
rect 20041 15039 20099 15045
rect 20257 15045 20269 15079
rect 20303 15076 20315 15079
rect 20622 15076 20628 15088
rect 20303 15048 20628 15076
rect 20303 15045 20315 15048
rect 20257 15039 20315 15045
rect 17221 15011 17279 15017
rect 17221 14977 17233 15011
rect 17267 14977 17279 15011
rect 17221 14971 17279 14977
rect 17405 15011 17463 15017
rect 17405 14977 17417 15011
rect 17451 14977 17463 15011
rect 17405 14971 17463 14977
rect 18233 15011 18291 15017
rect 18233 14977 18245 15011
rect 18279 14977 18291 15011
rect 18233 14971 18291 14977
rect 19061 15011 19119 15017
rect 19061 14977 19073 15011
rect 19107 15008 19119 15011
rect 19334 15008 19340 15020
rect 19107 14980 19340 15008
rect 19107 14977 19119 14980
rect 19061 14971 19119 14977
rect 17420 14940 17448 14971
rect 17052 14912 17448 14940
rect 16669 14903 16727 14909
rect 18248 14872 18276 14971
rect 19334 14968 19340 14980
rect 19392 14968 19398 15020
rect 18322 14900 18328 14952
rect 18380 14940 18386 14952
rect 20272 14940 20300 15039
rect 20622 15036 20628 15048
rect 20680 15036 20686 15088
rect 21910 15036 21916 15088
rect 21968 15076 21974 15088
rect 23569 15079 23627 15085
rect 23569 15076 23581 15079
rect 21968 15048 23581 15076
rect 21968 15036 21974 15048
rect 23569 15045 23581 15048
rect 23615 15076 23627 15079
rect 23934 15076 23940 15088
rect 23615 15048 23940 15076
rect 23615 15045 23627 15048
rect 23569 15039 23627 15045
rect 23934 15036 23940 15048
rect 23992 15036 23998 15088
rect 24854 15076 24860 15088
rect 24815 15048 24860 15076
rect 24854 15036 24860 15048
rect 24912 15036 24918 15088
rect 20714 14968 20720 15020
rect 20772 15008 20778 15020
rect 20901 15011 20959 15017
rect 20772 14980 20817 15008
rect 20772 14968 20778 14980
rect 20901 14977 20913 15011
rect 20947 15008 20959 15011
rect 20990 15008 20996 15020
rect 20947 14980 20996 15008
rect 20947 14977 20959 14980
rect 20901 14971 20959 14977
rect 20990 14968 20996 14980
rect 21048 14968 21054 15020
rect 21174 14968 21180 15020
rect 21232 15008 21238 15020
rect 21361 15011 21419 15017
rect 21361 15008 21373 15011
rect 21232 14980 21373 15008
rect 21232 14968 21238 14980
rect 21361 14977 21373 14980
rect 21407 14977 21419 15011
rect 21361 14971 21419 14977
rect 21726 14968 21732 15020
rect 21784 15008 21790 15020
rect 21821 15011 21879 15017
rect 21821 15008 21833 15011
rect 21784 14980 21833 15008
rect 21784 14968 21790 14980
rect 21821 14977 21833 14980
rect 21867 14977 21879 15011
rect 21821 14971 21879 14977
rect 22557 15011 22615 15017
rect 22557 14977 22569 15011
rect 22603 15008 22615 15011
rect 23014 15008 23020 15020
rect 22603 14980 23020 15008
rect 22603 14977 22615 14980
rect 22557 14971 22615 14977
rect 23014 14968 23020 14980
rect 23072 14968 23078 15020
rect 23750 15008 23756 15020
rect 23311 14980 23756 15008
rect 20530 14940 20536 14952
rect 18380 14912 20300 14940
rect 20491 14912 20536 14940
rect 18380 14900 18386 14912
rect 20530 14900 20536 14912
rect 20588 14900 20594 14952
rect 22002 14940 22008 14952
rect 21915 14912 22008 14940
rect 22002 14900 22008 14912
rect 22060 14940 22066 14952
rect 22281 14943 22339 14949
rect 22281 14940 22293 14943
rect 22060 14912 22293 14940
rect 22060 14900 22066 14912
rect 22281 14909 22293 14912
rect 22327 14909 22339 14943
rect 22281 14903 22339 14909
rect 22922 14900 22928 14952
rect 22980 14940 22986 14952
rect 23311 14940 23339 14980
rect 23750 14968 23756 14980
rect 23808 14968 23814 15020
rect 22980 14912 23339 14940
rect 23385 14943 23443 14949
rect 22980 14900 22986 14912
rect 23385 14909 23397 14943
rect 23431 14940 23443 14943
rect 23566 14940 23572 14952
rect 23431 14912 23572 14940
rect 23431 14909 23443 14912
rect 23385 14903 23443 14909
rect 23566 14900 23572 14912
rect 23624 14900 23630 14952
rect 18782 14872 18788 14884
rect 16316 14844 18788 14872
rect 14292 14776 14688 14804
rect 14737 14807 14795 14813
rect 14737 14773 14749 14807
rect 14783 14804 14795 14807
rect 16040 14804 16068 14844
rect 18782 14832 18788 14844
rect 18840 14832 18846 14884
rect 19058 14832 19064 14884
rect 19116 14872 19122 14884
rect 19613 14875 19671 14881
rect 19116 14844 19564 14872
rect 19116 14832 19122 14844
rect 14783 14776 16068 14804
rect 14783 14773 14795 14776
rect 14737 14767 14795 14773
rect 17678 14764 17684 14816
rect 17736 14804 17742 14816
rect 17957 14807 18015 14813
rect 17957 14804 17969 14807
rect 17736 14776 17969 14804
rect 17736 14764 17742 14776
rect 17957 14773 17969 14776
rect 18003 14804 18015 14807
rect 18046 14804 18052 14816
rect 18003 14776 18052 14804
rect 18003 14773 18015 14776
rect 17957 14767 18015 14773
rect 18046 14764 18052 14776
rect 18104 14764 18110 14816
rect 18506 14804 18512 14816
rect 18467 14776 18512 14804
rect 18506 14764 18512 14776
rect 18564 14764 18570 14816
rect 18966 14764 18972 14816
rect 19024 14804 19030 14816
rect 19429 14807 19487 14813
rect 19429 14804 19441 14807
rect 19024 14776 19441 14804
rect 19024 14764 19030 14776
rect 19429 14773 19441 14776
rect 19475 14773 19487 14807
rect 19536 14804 19564 14844
rect 19613 14841 19625 14875
rect 19659 14872 19671 14875
rect 21082 14872 21088 14884
rect 19659 14844 21088 14872
rect 19659 14841 19671 14844
rect 19613 14835 19671 14841
rect 21082 14832 21088 14844
rect 21140 14832 21146 14884
rect 21174 14832 21180 14884
rect 21232 14872 21238 14884
rect 22020 14872 22048 14900
rect 24397 14875 24455 14881
rect 24397 14872 24409 14875
rect 21232 14844 22048 14872
rect 23216 14844 24409 14872
rect 21232 14832 21238 14844
rect 20073 14807 20131 14813
rect 20073 14804 20085 14807
rect 19536 14776 20085 14804
rect 19429 14767 19487 14773
rect 20073 14773 20085 14776
rect 20119 14804 20131 14807
rect 23216 14804 23244 14844
rect 24397 14841 24409 14844
rect 24443 14841 24455 14875
rect 24397 14835 24455 14841
rect 24026 14804 24032 14816
rect 20119 14776 23244 14804
rect 23987 14776 24032 14804
rect 20119 14773 20131 14776
rect 20073 14767 20131 14773
rect 24026 14764 24032 14776
rect 24084 14764 24090 14816
rect 1104 14714 28888 14736
rect 1104 14662 5582 14714
rect 5634 14662 5646 14714
rect 5698 14662 5710 14714
rect 5762 14662 5774 14714
rect 5826 14662 5838 14714
rect 5890 14662 14846 14714
rect 14898 14662 14910 14714
rect 14962 14662 14974 14714
rect 15026 14662 15038 14714
rect 15090 14662 15102 14714
rect 15154 14662 24110 14714
rect 24162 14662 24174 14714
rect 24226 14662 24238 14714
rect 24290 14662 24302 14714
rect 24354 14662 24366 14714
rect 24418 14662 28888 14714
rect 1104 14640 28888 14662
rect 11974 14560 11980 14612
rect 12032 14600 12038 14612
rect 12894 14600 12900 14612
rect 12032 14572 12900 14600
rect 12032 14560 12038 14572
rect 12894 14560 12900 14572
rect 12952 14560 12958 14612
rect 13078 14560 13084 14612
rect 13136 14600 13142 14612
rect 15105 14603 15163 14609
rect 13136 14572 14688 14600
rect 13136 14560 13142 14572
rect 7929 14535 7987 14541
rect 7929 14501 7941 14535
rect 7975 14532 7987 14535
rect 8662 14532 8668 14544
rect 7975 14504 8668 14532
rect 7975 14501 7987 14504
rect 7929 14495 7987 14501
rect 8662 14492 8668 14504
rect 8720 14492 8726 14544
rect 12618 14492 12624 14544
rect 12676 14532 12682 14544
rect 13538 14532 13544 14544
rect 12676 14504 13544 14532
rect 12676 14492 12682 14504
rect 13538 14492 13544 14504
rect 13596 14532 13602 14544
rect 13633 14535 13691 14541
rect 13633 14532 13645 14535
rect 13596 14504 13645 14532
rect 13596 14492 13602 14504
rect 13633 14501 13645 14504
rect 13679 14501 13691 14535
rect 14660 14532 14688 14572
rect 15105 14569 15117 14603
rect 15151 14600 15163 14603
rect 15470 14600 15476 14612
rect 15151 14572 15476 14600
rect 15151 14569 15163 14572
rect 15105 14563 15163 14569
rect 15470 14560 15476 14572
rect 15528 14560 15534 14612
rect 15562 14560 15568 14612
rect 15620 14600 15626 14612
rect 16025 14603 16083 14609
rect 15620 14572 15976 14600
rect 15620 14560 15626 14572
rect 15654 14532 15660 14544
rect 14660 14504 15660 14532
rect 13633 14495 13691 14501
rect 15488 14476 15516 14504
rect 15654 14492 15660 14504
rect 15712 14492 15718 14544
rect 15948 14532 15976 14572
rect 16025 14569 16037 14603
rect 16071 14600 16083 14603
rect 16758 14600 16764 14612
rect 16071 14572 16764 14600
rect 16071 14569 16083 14572
rect 16025 14563 16083 14569
rect 16758 14560 16764 14572
rect 16816 14560 16822 14612
rect 18046 14560 18052 14612
rect 18104 14600 18110 14612
rect 18874 14600 18880 14612
rect 18104 14572 18880 14600
rect 18104 14560 18110 14572
rect 18874 14560 18880 14572
rect 18932 14560 18938 14612
rect 19429 14603 19487 14609
rect 19429 14569 19441 14603
rect 19475 14600 19487 14603
rect 19518 14600 19524 14612
rect 19475 14572 19524 14600
rect 19475 14569 19487 14572
rect 19429 14563 19487 14569
rect 19518 14560 19524 14572
rect 19576 14560 19582 14612
rect 19613 14603 19671 14609
rect 19613 14569 19625 14603
rect 19659 14600 19671 14603
rect 19978 14600 19984 14612
rect 19659 14572 19984 14600
rect 19659 14569 19671 14572
rect 19613 14563 19671 14569
rect 19978 14560 19984 14572
rect 20036 14560 20042 14612
rect 21358 14600 21364 14612
rect 21319 14572 21364 14600
rect 21358 14560 21364 14572
rect 21416 14560 21422 14612
rect 22554 14600 22560 14612
rect 22515 14572 22560 14600
rect 22554 14560 22560 14572
rect 22612 14560 22618 14612
rect 23017 14603 23075 14609
rect 23017 14569 23029 14603
rect 23063 14600 23075 14603
rect 23106 14600 23112 14612
rect 23063 14572 23112 14600
rect 23063 14569 23075 14572
rect 23017 14563 23075 14569
rect 23106 14560 23112 14572
rect 23164 14560 23170 14612
rect 23474 14560 23480 14612
rect 23532 14600 23538 14612
rect 26050 14600 26056 14612
rect 23532 14572 26056 14600
rect 23532 14560 23538 14572
rect 26050 14560 26056 14572
rect 26108 14560 26114 14612
rect 16390 14532 16396 14544
rect 15948 14504 16396 14532
rect 16390 14492 16396 14504
rect 16448 14492 16454 14544
rect 16482 14492 16488 14544
rect 16540 14532 16546 14544
rect 16853 14535 16911 14541
rect 16853 14532 16865 14535
rect 16540 14504 16865 14532
rect 16540 14492 16546 14504
rect 16853 14501 16865 14504
rect 16899 14501 16911 14535
rect 16853 14495 16911 14501
rect 17770 14492 17776 14544
rect 17828 14532 17834 14544
rect 18598 14532 18604 14544
rect 17828 14504 18604 14532
rect 17828 14492 17834 14504
rect 18598 14492 18604 14504
rect 18656 14492 18662 14544
rect 18782 14532 18788 14544
rect 18743 14504 18788 14532
rect 18782 14492 18788 14504
rect 18840 14532 18846 14544
rect 20530 14532 20536 14544
rect 18840 14504 20536 14532
rect 18840 14492 18846 14504
rect 14093 14467 14151 14473
rect 14093 14464 14105 14467
rect 12406 14436 14105 14464
rect 4430 14356 4436 14408
rect 4488 14396 4494 14408
rect 6549 14399 6607 14405
rect 6549 14396 6561 14399
rect 4488 14368 6561 14396
rect 4488 14356 4494 14368
rect 6549 14365 6561 14368
rect 6595 14396 6607 14399
rect 8294 14396 8300 14408
rect 6595 14368 8300 14396
rect 6595 14365 6607 14368
rect 6549 14359 6607 14365
rect 8294 14356 8300 14368
rect 8352 14356 8358 14408
rect 9125 14399 9183 14405
rect 9125 14365 9137 14399
rect 9171 14396 9183 14399
rect 9398 14396 9404 14408
rect 9171 14368 9404 14396
rect 9171 14365 9183 14368
rect 9125 14359 9183 14365
rect 9398 14356 9404 14368
rect 9456 14356 9462 14408
rect 11333 14399 11391 14405
rect 11333 14365 11345 14399
rect 11379 14396 11391 14399
rect 11974 14396 11980 14408
rect 11379 14368 11980 14396
rect 11379 14365 11391 14368
rect 11333 14359 11391 14365
rect 11974 14356 11980 14368
rect 12032 14356 12038 14408
rect 6816 14331 6874 14337
rect 6816 14297 6828 14331
rect 6862 14328 6874 14331
rect 6914 14328 6920 14340
rect 6862 14300 6920 14328
rect 6862 14297 6874 14300
rect 6816 14291 6874 14297
rect 6914 14288 6920 14300
rect 6972 14288 6978 14340
rect 11600 14331 11658 14337
rect 11600 14297 11612 14331
rect 11646 14328 11658 14331
rect 12406 14328 12434 14436
rect 14093 14433 14105 14436
rect 14139 14433 14151 14467
rect 14093 14427 14151 14433
rect 14182 14424 14188 14476
rect 14240 14464 14246 14476
rect 14240 14436 14596 14464
rect 14240 14424 14246 14436
rect 13265 14399 13323 14405
rect 13265 14396 13277 14399
rect 11646 14300 12434 14328
rect 12728 14368 13277 14396
rect 11646 14297 11658 14300
rect 11600 14291 11658 14297
rect 8478 14220 8484 14272
rect 8536 14260 8542 14272
rect 9033 14263 9091 14269
rect 9033 14260 9045 14263
rect 8536 14232 9045 14260
rect 8536 14220 8542 14232
rect 9033 14229 9045 14232
rect 9079 14229 9091 14263
rect 9490 14260 9496 14272
rect 9451 14232 9496 14260
rect 9033 14223 9091 14229
rect 9490 14220 9496 14232
rect 9548 14220 9554 14272
rect 12728 14269 12756 14368
rect 13265 14365 13277 14368
rect 13311 14396 13323 14399
rect 13541 14399 13599 14405
rect 13541 14396 13553 14399
rect 13311 14368 13553 14396
rect 13311 14365 13323 14368
rect 13265 14359 13323 14365
rect 13541 14365 13553 14368
rect 13587 14365 13599 14399
rect 13541 14359 13599 14365
rect 14274 14356 14280 14408
rect 14332 14396 14338 14408
rect 14568 14405 14596 14436
rect 15470 14424 15476 14476
rect 15528 14424 15534 14476
rect 15933 14467 15991 14473
rect 15933 14433 15945 14467
rect 15979 14464 15991 14467
rect 16022 14464 16028 14476
rect 15979 14436 16028 14464
rect 15979 14433 15991 14436
rect 15933 14427 15991 14433
rect 16022 14424 16028 14436
rect 16080 14424 16086 14476
rect 16114 14424 16120 14476
rect 16172 14464 16178 14476
rect 16172 14436 16217 14464
rect 16172 14424 16178 14436
rect 14369 14399 14427 14405
rect 14369 14396 14381 14399
rect 14332 14368 14381 14396
rect 14332 14356 14338 14368
rect 14369 14365 14381 14368
rect 14415 14365 14427 14399
rect 14369 14359 14427 14365
rect 14461 14399 14519 14405
rect 14461 14365 14473 14399
rect 14507 14365 14519 14399
rect 14461 14359 14519 14365
rect 14553 14399 14611 14405
rect 14553 14365 14565 14399
rect 14599 14365 14611 14399
rect 14553 14359 14611 14365
rect 14476 14328 14504 14359
rect 14642 14356 14648 14408
rect 14700 14396 14706 14408
rect 14737 14399 14795 14405
rect 14737 14396 14749 14399
rect 14700 14368 14749 14396
rect 14700 14356 14706 14368
rect 14737 14365 14749 14368
rect 14783 14365 14795 14399
rect 14737 14359 14795 14365
rect 15289 14399 15347 14405
rect 15289 14365 15301 14399
rect 15335 14396 15347 14399
rect 15378 14396 15384 14408
rect 15335 14368 15384 14396
rect 15335 14365 15347 14368
rect 15289 14359 15347 14365
rect 15378 14356 15384 14368
rect 15436 14396 15442 14408
rect 16301 14399 16359 14405
rect 15436 14368 15976 14396
rect 15436 14356 15442 14368
rect 15948 14340 15976 14368
rect 16301 14365 16313 14399
rect 16347 14396 16359 14399
rect 16500 14396 16528 14492
rect 18322 14464 18328 14476
rect 16960 14436 18328 14464
rect 16960 14408 16988 14436
rect 18322 14424 18328 14436
rect 18380 14424 18386 14476
rect 19334 14464 19340 14476
rect 19295 14436 19340 14464
rect 19334 14424 19340 14436
rect 19392 14424 19398 14476
rect 19996 14473 20024 14504
rect 20530 14492 20536 14504
rect 20588 14492 20594 14544
rect 20622 14492 20628 14544
rect 20680 14532 20686 14544
rect 24026 14532 24032 14544
rect 20680 14504 24032 14532
rect 20680 14492 20686 14504
rect 24026 14492 24032 14504
rect 24084 14492 24090 14544
rect 19981 14467 20039 14473
rect 19981 14433 19993 14467
rect 20027 14433 20039 14467
rect 19981 14427 20039 14433
rect 21450 14424 21456 14476
rect 21508 14464 21514 14476
rect 22189 14467 22247 14473
rect 21508 14436 22140 14464
rect 21508 14424 21514 14436
rect 16347 14368 16528 14396
rect 16761 14399 16819 14405
rect 16347 14365 16359 14368
rect 16301 14359 16359 14365
rect 16761 14365 16773 14399
rect 16807 14365 16819 14399
rect 16942 14396 16948 14408
rect 16855 14368 16948 14396
rect 16761 14359 16819 14365
rect 15194 14328 15200 14340
rect 14476 14300 15200 14328
rect 15194 14288 15200 14300
rect 15252 14288 15258 14340
rect 15473 14331 15531 14337
rect 15473 14297 15485 14331
rect 15519 14297 15531 14331
rect 15473 14291 15531 14297
rect 12713 14263 12771 14269
rect 12713 14229 12725 14263
rect 12759 14229 12771 14263
rect 12713 14223 12771 14229
rect 13906 14220 13912 14272
rect 13964 14260 13970 14272
rect 14274 14260 14280 14272
rect 13964 14232 14280 14260
rect 13964 14220 13970 14232
rect 14274 14220 14280 14232
rect 14332 14220 14338 14272
rect 14458 14220 14464 14272
rect 14516 14260 14522 14272
rect 14642 14260 14648 14272
rect 14516 14232 14648 14260
rect 14516 14220 14522 14232
rect 14642 14220 14648 14232
rect 14700 14220 14706 14272
rect 15488 14260 15516 14291
rect 15930 14288 15936 14340
rect 15988 14288 15994 14340
rect 16390 14288 16396 14340
rect 16448 14328 16454 14340
rect 16776 14328 16804 14359
rect 16942 14356 16948 14368
rect 17000 14356 17006 14408
rect 17034 14356 17040 14408
rect 17092 14396 17098 14408
rect 17681 14399 17739 14405
rect 17681 14396 17693 14399
rect 17092 14368 17693 14396
rect 17092 14356 17098 14368
rect 17681 14365 17693 14368
rect 17727 14396 17739 14399
rect 17862 14396 17868 14408
rect 17727 14368 17868 14396
rect 17727 14365 17739 14368
rect 17681 14359 17739 14365
rect 17862 14356 17868 14368
rect 17920 14356 17926 14408
rect 18046 14396 18052 14408
rect 18007 14368 18052 14396
rect 18046 14356 18052 14368
rect 18104 14356 18110 14408
rect 18166 14399 18224 14405
rect 18166 14365 18178 14399
rect 18212 14396 18224 14399
rect 18506 14396 18512 14408
rect 18212 14368 18512 14396
rect 18212 14365 18224 14368
rect 18166 14359 18224 14365
rect 18506 14356 18512 14368
rect 18564 14396 18570 14408
rect 18601 14399 18659 14405
rect 18601 14396 18613 14399
rect 18564 14368 18613 14396
rect 18564 14356 18570 14368
rect 18601 14365 18613 14368
rect 18647 14365 18659 14399
rect 19242 14396 19248 14408
rect 19203 14368 19248 14396
rect 18601 14359 18659 14365
rect 19242 14356 19248 14368
rect 19300 14356 19306 14408
rect 20162 14396 20168 14408
rect 20123 14368 20168 14396
rect 20162 14356 20168 14368
rect 20220 14396 20226 14408
rect 20625 14399 20683 14405
rect 20625 14396 20637 14399
rect 20220 14368 20637 14396
rect 20220 14356 20226 14368
rect 20625 14365 20637 14368
rect 20671 14365 20683 14399
rect 21174 14396 21180 14408
rect 21135 14368 21180 14396
rect 20625 14359 20683 14365
rect 21174 14356 21180 14368
rect 21232 14356 21238 14408
rect 21634 14356 21640 14408
rect 21692 14396 21698 14408
rect 21821 14399 21879 14405
rect 21821 14396 21833 14399
rect 21692 14368 21833 14396
rect 21692 14356 21698 14368
rect 21821 14365 21833 14368
rect 21867 14365 21879 14399
rect 22002 14396 22008 14408
rect 21963 14368 22008 14396
rect 21821 14359 21879 14365
rect 22002 14356 22008 14368
rect 22060 14356 22066 14408
rect 22112 14396 22140 14436
rect 22189 14433 22201 14467
rect 22235 14464 22247 14467
rect 22235 14436 23612 14464
rect 22235 14433 22247 14436
rect 22189 14427 22247 14433
rect 22465 14399 22523 14405
rect 22465 14396 22477 14399
rect 22112 14368 22477 14396
rect 22465 14365 22477 14368
rect 22511 14365 22523 14399
rect 22646 14396 22652 14408
rect 22607 14368 22652 14396
rect 22465 14359 22523 14365
rect 22646 14356 22652 14368
rect 22704 14396 22710 14408
rect 23584 14405 23612 14436
rect 22925 14399 22983 14405
rect 22925 14396 22937 14399
rect 22704 14368 22937 14396
rect 22704 14356 22710 14368
rect 22925 14365 22937 14368
rect 22971 14365 22983 14399
rect 22925 14359 22983 14365
rect 23109 14399 23167 14405
rect 23109 14365 23121 14399
rect 23155 14365 23167 14399
rect 23109 14359 23167 14365
rect 23569 14399 23627 14405
rect 23569 14365 23581 14399
rect 23615 14365 23627 14399
rect 23842 14396 23848 14408
rect 23803 14368 23848 14396
rect 23569 14359 23627 14365
rect 17957 14331 18015 14337
rect 17957 14328 17969 14331
rect 16448 14300 17969 14328
rect 16448 14288 16454 14300
rect 17957 14297 17969 14300
rect 18003 14328 18015 14331
rect 19058 14328 19064 14340
rect 18003 14300 19064 14328
rect 18003 14297 18015 14300
rect 17957 14291 18015 14297
rect 19058 14288 19064 14300
rect 19116 14288 19122 14340
rect 20180 14300 20484 14328
rect 15746 14260 15752 14272
rect 15488 14232 15752 14260
rect 15746 14220 15752 14232
rect 15804 14260 15810 14272
rect 16209 14263 16267 14269
rect 16209 14260 16221 14263
rect 15804 14232 16221 14260
rect 15804 14220 15810 14232
rect 16209 14229 16221 14232
rect 16255 14229 16267 14263
rect 16209 14223 16267 14229
rect 18325 14263 18383 14269
rect 18325 14229 18337 14263
rect 18371 14260 18383 14263
rect 18414 14260 18420 14272
rect 18371 14232 18420 14260
rect 18371 14229 18383 14232
rect 18325 14223 18383 14229
rect 18414 14220 18420 14232
rect 18472 14220 18478 14272
rect 18874 14220 18880 14272
rect 18932 14260 18938 14272
rect 20180 14260 20208 14300
rect 20346 14260 20352 14272
rect 18932 14232 20208 14260
rect 20307 14232 20352 14260
rect 18932 14220 18938 14232
rect 20346 14220 20352 14232
rect 20404 14220 20410 14272
rect 20456 14260 20484 14300
rect 20530 14288 20536 14340
rect 20588 14328 20594 14340
rect 20809 14331 20867 14337
rect 20809 14328 20821 14331
rect 20588 14300 20821 14328
rect 20588 14288 20594 14300
rect 20809 14297 20821 14300
rect 20855 14297 20867 14331
rect 20809 14291 20867 14297
rect 20990 14288 20996 14340
rect 21048 14328 21054 14340
rect 22370 14328 22376 14340
rect 21048 14300 22376 14328
rect 21048 14288 21054 14300
rect 22370 14288 22376 14300
rect 22428 14328 22434 14340
rect 23124 14328 23152 14359
rect 23842 14356 23848 14368
rect 23900 14356 23906 14408
rect 23934 14356 23940 14408
rect 23992 14396 23998 14408
rect 25777 14399 25835 14405
rect 25777 14396 25789 14399
rect 23992 14368 25789 14396
rect 23992 14356 23998 14368
rect 25777 14365 25789 14368
rect 25823 14396 25835 14399
rect 26053 14399 26111 14405
rect 26053 14396 26065 14399
rect 25823 14368 26065 14396
rect 25823 14365 25835 14368
rect 25777 14359 25835 14365
rect 26053 14365 26065 14368
rect 26099 14365 26111 14399
rect 26053 14359 26111 14365
rect 25510 14331 25568 14337
rect 25510 14328 25522 14331
rect 22428 14300 23152 14328
rect 24044 14300 25522 14328
rect 22428 14288 22434 14300
rect 20714 14260 20720 14272
rect 20456 14232 20720 14260
rect 20714 14220 20720 14232
rect 20772 14220 20778 14272
rect 23382 14260 23388 14272
rect 23343 14232 23388 14260
rect 23382 14220 23388 14232
rect 23440 14220 23446 14272
rect 24044 14269 24072 14300
rect 25510 14297 25522 14300
rect 25556 14297 25568 14331
rect 25510 14291 25568 14297
rect 25866 14288 25872 14340
rect 25924 14328 25930 14340
rect 26298 14331 26356 14337
rect 26298 14328 26310 14331
rect 25924 14300 26310 14328
rect 25924 14288 25930 14300
rect 26298 14297 26310 14300
rect 26344 14297 26356 14331
rect 26298 14291 26356 14297
rect 24029 14263 24087 14269
rect 24029 14229 24041 14263
rect 24075 14229 24087 14263
rect 24029 14223 24087 14229
rect 24397 14263 24455 14269
rect 24397 14229 24409 14263
rect 24443 14260 24455 14263
rect 24486 14260 24492 14272
rect 24443 14232 24492 14260
rect 24443 14229 24455 14232
rect 24397 14223 24455 14229
rect 24486 14220 24492 14232
rect 24544 14220 24550 14272
rect 27433 14263 27491 14269
rect 27433 14229 27445 14263
rect 27479 14260 27491 14263
rect 28074 14260 28080 14272
rect 27479 14232 28080 14260
rect 27479 14229 27491 14232
rect 27433 14223 27491 14229
rect 28074 14220 28080 14232
rect 28132 14220 28138 14272
rect 1104 14170 28888 14192
rect 1104 14118 10214 14170
rect 10266 14118 10278 14170
rect 10330 14118 10342 14170
rect 10394 14118 10406 14170
rect 10458 14118 10470 14170
rect 10522 14118 19478 14170
rect 19530 14118 19542 14170
rect 19594 14118 19606 14170
rect 19658 14118 19670 14170
rect 19722 14118 19734 14170
rect 19786 14118 28888 14170
rect 1104 14096 28888 14118
rect 6914 14016 6920 14068
rect 6972 14056 6978 14068
rect 6972 14028 7017 14056
rect 6972 14016 6978 14028
rect 8110 14016 8116 14068
rect 8168 14056 8174 14068
rect 8205 14059 8263 14065
rect 8205 14056 8217 14059
rect 8168 14028 8217 14056
rect 8168 14016 8174 14028
rect 8205 14025 8217 14028
rect 8251 14025 8263 14059
rect 13078 14056 13084 14068
rect 8205 14019 8263 14025
rect 12268 14028 13084 14056
rect 6546 13948 6552 14000
rect 6604 13988 6610 14000
rect 6641 13991 6699 13997
rect 6641 13988 6653 13991
rect 6604 13960 6653 13988
rect 6604 13948 6610 13960
rect 6641 13957 6653 13960
rect 6687 13988 6699 13991
rect 6687 13960 7880 13988
rect 6687 13957 6699 13960
rect 6641 13951 6699 13957
rect 4884 13923 4942 13929
rect 4884 13889 4896 13923
rect 4930 13920 4942 13923
rect 6270 13920 6276 13932
rect 4930 13892 6276 13920
rect 4930 13889 4942 13892
rect 4884 13883 4942 13889
rect 6270 13880 6276 13892
rect 6328 13880 6334 13932
rect 7098 13920 7104 13932
rect 7059 13892 7104 13920
rect 7098 13880 7104 13892
rect 7156 13880 7162 13932
rect 7561 13923 7619 13929
rect 7561 13889 7573 13923
rect 7607 13889 7619 13923
rect 7852 13920 7880 13960
rect 8018 13948 8024 14000
rect 8076 13988 8082 14000
rect 9125 13991 9183 13997
rect 9125 13988 9137 13991
rect 8076 13960 9137 13988
rect 8076 13948 8082 13960
rect 9125 13957 9137 13960
rect 9171 13957 9183 13991
rect 10134 13988 10140 14000
rect 9125 13951 9183 13957
rect 9232 13960 10140 13988
rect 8478 13920 8484 13932
rect 7852 13892 8248 13920
rect 8439 13892 8484 13920
rect 7561 13883 7619 13889
rect 1394 13852 1400 13864
rect 1355 13824 1400 13852
rect 1394 13812 1400 13824
rect 1452 13812 1458 13864
rect 4430 13812 4436 13864
rect 4488 13852 4494 13864
rect 4617 13855 4675 13861
rect 4617 13852 4629 13855
rect 4488 13824 4629 13852
rect 4488 13812 4494 13824
rect 4617 13821 4629 13824
rect 4663 13821 4675 13855
rect 4617 13815 4675 13821
rect 6730 13812 6736 13864
rect 6788 13852 6794 13864
rect 7469 13855 7527 13861
rect 7469 13852 7481 13855
rect 6788 13824 7481 13852
rect 6788 13812 6794 13824
rect 7469 13821 7481 13824
rect 7515 13821 7527 13855
rect 7469 13815 7527 13821
rect 7576 13852 7604 13883
rect 8110 13852 8116 13864
rect 7576 13824 8116 13852
rect 5997 13787 6055 13793
rect 5997 13753 6009 13787
rect 6043 13784 6055 13787
rect 6043 13756 6684 13784
rect 6043 13753 6055 13756
rect 5997 13747 6055 13753
rect 6656 13716 6684 13756
rect 7006 13716 7012 13728
rect 6656 13688 7012 13716
rect 7006 13676 7012 13688
rect 7064 13716 7070 13728
rect 7576 13716 7604 13824
rect 8110 13812 8116 13824
rect 8168 13812 8174 13864
rect 8220 13784 8248 13892
rect 8478 13880 8484 13892
rect 8536 13880 8542 13932
rect 8570 13880 8576 13932
rect 8628 13920 8634 13932
rect 8938 13920 8944 13932
rect 8628 13892 8673 13920
rect 8899 13892 8944 13920
rect 8628 13880 8634 13892
rect 8938 13880 8944 13892
rect 8996 13880 9002 13932
rect 9232 13929 9260 13960
rect 10134 13948 10140 13960
rect 10192 13948 10198 14000
rect 9217 13923 9275 13929
rect 9217 13889 9229 13923
rect 9263 13889 9275 13923
rect 9217 13883 9275 13889
rect 9582 13880 9588 13932
rect 9640 13920 9646 13932
rect 9749 13923 9807 13929
rect 9749 13920 9761 13923
rect 9640 13892 9761 13920
rect 9640 13880 9646 13892
rect 9749 13889 9761 13892
rect 9795 13889 9807 13923
rect 11698 13920 11704 13932
rect 11659 13892 11704 13920
rect 9749 13883 9807 13889
rect 11698 13880 11704 13892
rect 11756 13880 11762 13932
rect 12158 13920 12164 13932
rect 12119 13892 12164 13920
rect 12158 13880 12164 13892
rect 12216 13880 12222 13932
rect 12268 13929 12296 14028
rect 13078 14016 13084 14028
rect 13136 14016 13142 14068
rect 13170 14016 13176 14068
rect 13228 14056 13234 14068
rect 13228 14028 13273 14056
rect 13464 14028 13952 14056
rect 13228 14016 13234 14028
rect 12434 13948 12440 14000
rect 12492 13988 12498 14000
rect 13464 13997 13492 14028
rect 13449 13991 13507 13997
rect 12492 13960 12537 13988
rect 12492 13948 12498 13960
rect 13449 13957 13461 13991
rect 13495 13957 13507 13991
rect 13924 13988 13952 14028
rect 15194 14016 15200 14068
rect 15252 14056 15258 14068
rect 15378 14056 15384 14068
rect 15252 14028 15384 14056
rect 15252 14016 15258 14028
rect 15378 14016 15384 14028
rect 15436 14056 15442 14068
rect 16209 14059 16267 14065
rect 16209 14056 16221 14059
rect 15436 14028 16221 14056
rect 15436 14016 15442 14028
rect 16209 14025 16221 14028
rect 16255 14025 16267 14059
rect 18601 14059 18659 14065
rect 18601 14056 18613 14059
rect 16209 14019 16267 14025
rect 18156 14028 18613 14056
rect 14614 13991 14672 13997
rect 14614 13988 14626 13991
rect 13924 13960 14626 13988
rect 13449 13951 13507 13957
rect 14614 13957 14626 13960
rect 14660 13957 14672 13991
rect 14614 13951 14672 13957
rect 15838 13948 15844 14000
rect 15896 13988 15902 14000
rect 18156 13997 18184 14028
rect 18601 14025 18613 14028
rect 18647 14056 18659 14059
rect 19242 14056 19248 14068
rect 18647 14028 19248 14056
rect 18647 14025 18659 14028
rect 18601 14019 18659 14025
rect 19242 14016 19248 14028
rect 19300 14016 19306 14068
rect 20346 14016 20352 14068
rect 20404 14056 20410 14068
rect 25777 14059 25835 14065
rect 20404 14028 25636 14056
rect 20404 14016 20410 14028
rect 18141 13991 18199 13997
rect 15896 13960 18092 13988
rect 15896 13948 15902 13960
rect 12254 13923 12312 13929
rect 12254 13889 12266 13923
rect 12300 13889 12312 13923
rect 12526 13920 12532 13932
rect 12487 13892 12532 13920
rect 12254 13883 12312 13889
rect 12526 13880 12532 13892
rect 12584 13880 12590 13932
rect 12667 13923 12725 13929
rect 12667 13889 12679 13923
rect 12713 13920 12725 13923
rect 13354 13920 13360 13932
rect 12713 13892 13360 13920
rect 12713 13889 12725 13892
rect 12667 13883 12725 13889
rect 13354 13880 13360 13892
rect 13412 13880 13418 13932
rect 13722 13920 13728 13932
rect 13683 13892 13728 13920
rect 13722 13880 13728 13892
rect 13780 13880 13786 13932
rect 13817 13923 13875 13929
rect 13817 13889 13829 13923
rect 13863 13889 13875 13923
rect 13817 13883 13875 13889
rect 8294 13812 8300 13864
rect 8352 13852 8358 13864
rect 9493 13855 9551 13861
rect 9493 13852 9505 13855
rect 8352 13824 9505 13852
rect 8352 13812 8358 13824
rect 9493 13821 9505 13824
rect 9539 13821 9551 13855
rect 9493 13815 9551 13821
rect 11793 13787 11851 13793
rect 8220 13756 9536 13784
rect 8202 13716 8208 13728
rect 7064 13688 7604 13716
rect 8163 13688 8208 13716
rect 7064 13676 7070 13688
rect 8202 13676 8208 13688
rect 8260 13676 8266 13728
rect 8312 13725 8340 13756
rect 9508 13728 9536 13756
rect 11793 13753 11805 13787
rect 11839 13784 11851 13787
rect 12434 13784 12440 13796
rect 11839 13756 12440 13784
rect 11839 13753 11851 13756
rect 11793 13747 11851 13753
rect 12434 13744 12440 13756
rect 12492 13744 12498 13796
rect 13630 13744 13636 13796
rect 13688 13784 13694 13796
rect 13832 13784 13860 13883
rect 13906 13880 13912 13932
rect 13964 13920 13970 13932
rect 14093 13923 14151 13929
rect 13964 13892 14009 13920
rect 13964 13880 13970 13892
rect 14093 13889 14105 13923
rect 14139 13920 14151 13923
rect 14458 13920 14464 13932
rect 14139 13892 14464 13920
rect 14139 13889 14151 13892
rect 14093 13883 14151 13889
rect 14458 13880 14464 13892
rect 14516 13880 14522 13932
rect 15654 13880 15660 13932
rect 15712 13920 15718 13932
rect 16117 13923 16175 13929
rect 16117 13920 16129 13923
rect 15712 13892 16129 13920
rect 15712 13880 15718 13892
rect 16117 13889 16129 13892
rect 16163 13920 16175 13923
rect 16945 13923 17003 13929
rect 16945 13920 16957 13923
rect 16163 13892 16957 13920
rect 16163 13889 16175 13892
rect 16117 13883 16175 13889
rect 16945 13889 16957 13892
rect 16991 13889 17003 13923
rect 16945 13883 17003 13889
rect 17034 13880 17040 13932
rect 17092 13920 17098 13932
rect 17770 13920 17776 13932
rect 17092 13892 17776 13920
rect 17092 13880 17098 13892
rect 17770 13880 17776 13892
rect 17828 13880 17834 13932
rect 14369 13855 14427 13861
rect 14369 13852 14381 13855
rect 13688 13756 13860 13784
rect 13924 13824 14381 13852
rect 13688 13744 13694 13756
rect 8297 13719 8355 13725
rect 8297 13685 8309 13719
rect 8343 13685 8355 13719
rect 8297 13679 8355 13685
rect 8386 13676 8392 13728
rect 8444 13716 8450 13728
rect 9033 13719 9091 13725
rect 8444 13688 8489 13716
rect 8444 13676 8450 13688
rect 9033 13685 9045 13719
rect 9079 13716 9091 13719
rect 9122 13716 9128 13728
rect 9079 13688 9128 13716
rect 9079 13685 9091 13688
rect 9033 13679 9091 13685
rect 9122 13676 9128 13688
rect 9180 13676 9186 13728
rect 9490 13676 9496 13728
rect 9548 13676 9554 13728
rect 10226 13676 10232 13728
rect 10284 13716 10290 13728
rect 10873 13719 10931 13725
rect 10873 13716 10885 13719
rect 10284 13688 10885 13716
rect 10284 13676 10290 13688
rect 10873 13685 10885 13688
rect 10919 13716 10931 13719
rect 11698 13716 11704 13728
rect 10919 13688 11704 13716
rect 10919 13685 10931 13688
rect 10873 13679 10931 13685
rect 11698 13676 11704 13688
rect 11756 13676 11762 13728
rect 12802 13716 12808 13728
rect 12763 13688 12808 13716
rect 12802 13676 12808 13688
rect 12860 13676 12866 13728
rect 13722 13676 13728 13728
rect 13780 13716 13786 13728
rect 13924 13716 13952 13824
rect 14369 13821 14381 13824
rect 14415 13821 14427 13855
rect 16666 13852 16672 13864
rect 16627 13824 16672 13852
rect 14369 13815 14427 13821
rect 16666 13812 16672 13824
rect 16724 13812 16730 13864
rect 18064 13852 18092 13960
rect 18141 13957 18153 13991
rect 18187 13957 18199 13991
rect 18141 13951 18199 13957
rect 18322 13948 18328 14000
rect 18380 13988 18386 14000
rect 18380 13960 18644 13988
rect 18380 13948 18386 13960
rect 18414 13920 18420 13932
rect 18375 13892 18420 13920
rect 18414 13880 18420 13892
rect 18472 13880 18478 13932
rect 18616 13929 18644 13960
rect 18874 13948 18880 14000
rect 18932 13988 18938 14000
rect 19521 13991 19579 13997
rect 19521 13988 19533 13991
rect 18932 13960 19533 13988
rect 18932 13948 18938 13960
rect 19521 13957 19533 13960
rect 19567 13957 19579 13991
rect 19521 13951 19579 13957
rect 20073 13991 20131 13997
rect 20073 13957 20085 13991
rect 20119 13988 20131 13991
rect 20530 13988 20536 14000
rect 20119 13960 20536 13988
rect 20119 13957 20131 13960
rect 20073 13951 20131 13957
rect 20530 13948 20536 13960
rect 20588 13948 20594 14000
rect 22956 13991 23014 13997
rect 22956 13957 22968 13991
rect 23002 13988 23014 13991
rect 23382 13988 23388 14000
rect 23002 13960 23388 13988
rect 23002 13957 23014 13960
rect 22956 13951 23014 13957
rect 23382 13948 23388 13960
rect 23440 13948 23446 14000
rect 23492 13960 25084 13988
rect 18601 13923 18659 13929
rect 18601 13889 18613 13923
rect 18647 13920 18659 13923
rect 18969 13923 19027 13929
rect 18969 13920 18981 13923
rect 18647 13892 18981 13920
rect 18647 13889 18659 13892
rect 18601 13883 18659 13889
rect 18969 13889 18981 13892
rect 19015 13889 19027 13923
rect 18969 13883 19027 13889
rect 19978 13880 19984 13932
rect 20036 13920 20042 13932
rect 20625 13923 20683 13929
rect 20625 13920 20637 13923
rect 20036 13892 20637 13920
rect 20036 13880 20042 13892
rect 20625 13889 20637 13892
rect 20671 13889 20683 13923
rect 20898 13920 20904 13932
rect 20859 13892 20904 13920
rect 20625 13883 20683 13889
rect 20640 13852 20668 13883
rect 20898 13880 20904 13892
rect 20956 13880 20962 13932
rect 21085 13923 21143 13929
rect 21085 13889 21097 13923
rect 21131 13920 21143 13923
rect 21174 13920 21180 13932
rect 21131 13892 21180 13920
rect 21131 13889 21143 13892
rect 21085 13883 21143 13889
rect 21174 13880 21180 13892
rect 21232 13880 21238 13932
rect 23492 13920 23520 13960
rect 22066 13892 23520 13920
rect 22066 13852 22094 13892
rect 23566 13880 23572 13932
rect 23624 13920 23630 13932
rect 24029 13923 24087 13929
rect 24029 13920 24041 13923
rect 23624 13892 24041 13920
rect 23624 13880 23630 13892
rect 24029 13889 24041 13892
rect 24075 13889 24087 13923
rect 24029 13883 24087 13889
rect 24121 13923 24179 13929
rect 24121 13889 24133 13923
rect 24167 13920 24179 13923
rect 24486 13920 24492 13932
rect 24167 13892 24492 13920
rect 24167 13889 24179 13892
rect 24121 13883 24179 13889
rect 24486 13880 24492 13892
rect 24544 13880 24550 13932
rect 24946 13920 24952 13932
rect 24907 13892 24952 13920
rect 24946 13880 24952 13892
rect 25004 13880 25010 13932
rect 25056 13864 25084 13960
rect 25608 13929 25636 14028
rect 25777 14025 25789 14059
rect 25823 14056 25835 14059
rect 25866 14056 25872 14068
rect 25823 14028 25872 14056
rect 25823 14025 25835 14028
rect 25777 14019 25835 14025
rect 25866 14016 25872 14028
rect 25924 14016 25930 14068
rect 26050 14056 26056 14068
rect 26011 14028 26056 14056
rect 26050 14016 26056 14028
rect 26108 14016 26114 14068
rect 26418 14056 26424 14068
rect 26379 14028 26424 14056
rect 26418 14016 26424 14028
rect 26476 14016 26482 14068
rect 25593 13923 25651 13929
rect 25593 13889 25605 13923
rect 25639 13889 25651 13923
rect 25593 13883 25651 13889
rect 27801 13923 27859 13929
rect 27801 13889 27813 13923
rect 27847 13920 27859 13923
rect 28258 13920 28264 13932
rect 27847 13892 28264 13920
rect 27847 13889 27859 13892
rect 27801 13883 27859 13889
rect 28258 13880 28264 13892
rect 28316 13880 28322 13932
rect 18064 13824 19334 13852
rect 20640 13824 22094 13852
rect 23201 13855 23259 13861
rect 16022 13744 16028 13796
rect 16080 13784 16086 13796
rect 16390 13784 16396 13796
rect 16080 13756 16396 13784
rect 16080 13744 16086 13756
rect 16390 13744 16396 13756
rect 16448 13784 16454 13796
rect 17865 13787 17923 13793
rect 17865 13784 17877 13787
rect 16448 13756 17877 13784
rect 16448 13744 16454 13756
rect 17865 13753 17877 13756
rect 17911 13753 17923 13787
rect 17865 13747 17923 13753
rect 13780 13688 13952 13716
rect 13780 13676 13786 13688
rect 14182 13676 14188 13728
rect 14240 13716 14246 13728
rect 14642 13716 14648 13728
rect 14240 13688 14648 13716
rect 14240 13676 14246 13688
rect 14642 13676 14648 13688
rect 14700 13716 14706 13728
rect 15749 13719 15807 13725
rect 15749 13716 15761 13719
rect 14700 13688 15761 13716
rect 14700 13676 14706 13688
rect 15749 13685 15761 13688
rect 15795 13685 15807 13719
rect 17954 13716 17960 13728
rect 17915 13688 17960 13716
rect 15749 13679 15807 13685
rect 17954 13676 17960 13688
rect 18012 13676 18018 13728
rect 18138 13716 18144 13728
rect 18099 13688 18144 13716
rect 18138 13676 18144 13688
rect 18196 13676 18202 13728
rect 18598 13676 18604 13728
rect 18656 13716 18662 13728
rect 18969 13719 19027 13725
rect 18969 13716 18981 13719
rect 18656 13688 18981 13716
rect 18656 13676 18662 13688
rect 18969 13685 18981 13688
rect 19015 13685 19027 13719
rect 19306 13716 19334 13824
rect 23201 13821 23213 13855
rect 23247 13852 23259 13855
rect 23934 13852 23940 13864
rect 23247 13824 23940 13852
rect 23247 13821 23259 13824
rect 23201 13815 23259 13821
rect 23934 13812 23940 13824
rect 23992 13812 23998 13864
rect 24213 13855 24271 13861
rect 24213 13821 24225 13855
rect 24259 13821 24271 13855
rect 24213 13815 24271 13821
rect 23382 13744 23388 13796
rect 23440 13784 23446 13796
rect 24228 13784 24256 13815
rect 24670 13812 24676 13864
rect 24728 13852 24734 13864
rect 24765 13855 24823 13861
rect 24765 13852 24777 13855
rect 24728 13824 24777 13852
rect 24728 13812 24734 13824
rect 24765 13821 24777 13824
rect 24811 13821 24823 13855
rect 24765 13815 24823 13821
rect 25038 13812 25044 13864
rect 25096 13852 25102 13864
rect 28077 13855 28135 13861
rect 28077 13852 28089 13855
rect 25096 13824 28089 13852
rect 25096 13812 25102 13824
rect 28077 13821 28089 13824
rect 28123 13821 28135 13855
rect 28077 13815 28135 13821
rect 23440 13756 24256 13784
rect 23440 13744 23446 13756
rect 19981 13719 20039 13725
rect 19981 13716 19993 13719
rect 19306 13688 19993 13716
rect 18969 13679 19027 13685
rect 19981 13685 19993 13688
rect 20027 13716 20039 13719
rect 21726 13716 21732 13728
rect 20027 13688 21732 13716
rect 20027 13685 20039 13688
rect 19981 13679 20039 13685
rect 21726 13676 21732 13688
rect 21784 13676 21790 13728
rect 21821 13719 21879 13725
rect 21821 13685 21833 13719
rect 21867 13716 21879 13719
rect 22554 13716 22560 13728
rect 21867 13688 22560 13716
rect 21867 13685 21879 13688
rect 21821 13679 21879 13685
rect 22554 13676 22560 13688
rect 22612 13676 22618 13728
rect 23658 13716 23664 13728
rect 23619 13688 23664 13716
rect 23658 13676 23664 13688
rect 23716 13676 23722 13728
rect 25133 13719 25191 13725
rect 25133 13685 25145 13719
rect 25179 13716 25191 13719
rect 25406 13716 25412 13728
rect 25179 13688 25412 13716
rect 25179 13685 25191 13688
rect 25133 13679 25191 13685
rect 25406 13676 25412 13688
rect 25464 13676 25470 13728
rect 1104 13626 28888 13648
rect 1104 13574 5582 13626
rect 5634 13574 5646 13626
rect 5698 13574 5710 13626
rect 5762 13574 5774 13626
rect 5826 13574 5838 13626
rect 5890 13574 14846 13626
rect 14898 13574 14910 13626
rect 14962 13574 14974 13626
rect 15026 13574 15038 13626
rect 15090 13574 15102 13626
rect 15154 13574 24110 13626
rect 24162 13574 24174 13626
rect 24226 13574 24238 13626
rect 24290 13574 24302 13626
rect 24354 13574 24366 13626
rect 24418 13574 28888 13626
rect 1104 13552 28888 13574
rect 6270 13512 6276 13524
rect 6231 13484 6276 13512
rect 6270 13472 6276 13484
rect 6328 13472 6334 13524
rect 6546 13512 6552 13524
rect 6507 13484 6552 13512
rect 6546 13472 6552 13484
rect 6604 13472 6610 13524
rect 7098 13472 7104 13524
rect 7156 13512 7162 13524
rect 7193 13515 7251 13521
rect 7193 13512 7205 13515
rect 7156 13484 7205 13512
rect 7156 13472 7162 13484
rect 7193 13481 7205 13484
rect 7239 13481 7251 13515
rect 7193 13475 7251 13481
rect 7377 13515 7435 13521
rect 7377 13481 7389 13515
rect 7423 13512 7435 13515
rect 7926 13512 7932 13524
rect 7423 13484 7932 13512
rect 7423 13481 7435 13484
rect 7377 13475 7435 13481
rect 7926 13472 7932 13484
rect 7984 13472 7990 13524
rect 8110 13472 8116 13524
rect 8168 13512 8174 13524
rect 9582 13512 9588 13524
rect 8168 13484 9352 13512
rect 9543 13484 9588 13512
rect 8168 13472 8174 13484
rect 6457 13447 6515 13453
rect 6457 13413 6469 13447
rect 6503 13444 6515 13447
rect 7650 13444 7656 13456
rect 6503 13416 7656 13444
rect 6503 13413 6515 13416
rect 6457 13407 6515 13413
rect 7650 13404 7656 13416
rect 7708 13444 7714 13456
rect 8202 13444 8208 13456
rect 7708 13416 8208 13444
rect 7708 13404 7714 13416
rect 8202 13404 8208 13416
rect 8260 13404 8266 13456
rect 6641 13379 6699 13385
rect 6641 13345 6653 13379
rect 6687 13376 6699 13379
rect 6822 13376 6828 13388
rect 6687 13348 6828 13376
rect 6687 13345 6699 13348
rect 6641 13339 6699 13345
rect 6822 13336 6828 13348
rect 6880 13336 6886 13388
rect 8021 13379 8079 13385
rect 8021 13345 8033 13379
rect 8067 13376 8079 13379
rect 8386 13376 8392 13388
rect 8067 13348 8392 13376
rect 8067 13345 8079 13348
rect 8021 13339 8079 13345
rect 8386 13336 8392 13348
rect 8444 13376 8450 13388
rect 9324 13376 9352 13484
rect 9582 13472 9588 13484
rect 9640 13472 9646 13524
rect 10045 13515 10103 13521
rect 10045 13481 10057 13515
rect 10091 13481 10103 13515
rect 10045 13475 10103 13481
rect 11333 13515 11391 13521
rect 11333 13481 11345 13515
rect 11379 13512 11391 13515
rect 12158 13512 12164 13524
rect 11379 13484 12164 13512
rect 11379 13481 11391 13484
rect 11333 13475 11391 13481
rect 9490 13404 9496 13456
rect 9548 13444 9554 13456
rect 10060 13444 10088 13475
rect 12158 13472 12164 13484
rect 12216 13472 12222 13524
rect 13906 13472 13912 13524
rect 13964 13512 13970 13524
rect 14185 13515 14243 13521
rect 14185 13512 14197 13515
rect 13964 13484 14197 13512
rect 13964 13472 13970 13484
rect 14185 13481 14197 13484
rect 14231 13481 14243 13515
rect 14185 13475 14243 13481
rect 14274 13472 14280 13524
rect 14332 13512 14338 13524
rect 14921 13515 14979 13521
rect 14921 13512 14933 13515
rect 14332 13484 14933 13512
rect 14332 13472 14338 13484
rect 14921 13481 14933 13484
rect 14967 13512 14979 13515
rect 15194 13512 15200 13524
rect 14967 13484 15200 13512
rect 14967 13481 14979 13484
rect 14921 13475 14979 13481
rect 15194 13472 15200 13484
rect 15252 13472 15258 13524
rect 15473 13515 15531 13521
rect 15473 13481 15485 13515
rect 15519 13512 15531 13515
rect 15562 13512 15568 13524
rect 15519 13484 15568 13512
rect 15519 13481 15531 13484
rect 15473 13475 15531 13481
rect 15562 13472 15568 13484
rect 15620 13472 15626 13524
rect 16577 13515 16635 13521
rect 16577 13481 16589 13515
rect 16623 13512 16635 13515
rect 16758 13512 16764 13524
rect 16623 13484 16764 13512
rect 16623 13481 16635 13484
rect 16577 13475 16635 13481
rect 16758 13472 16764 13484
rect 16816 13472 16822 13524
rect 17954 13512 17960 13524
rect 17144 13484 17960 13512
rect 9548 13416 10088 13444
rect 11624 13416 13768 13444
rect 9548 13404 9554 13416
rect 10873 13379 10931 13385
rect 10873 13376 10885 13379
rect 8444 13348 9260 13376
rect 9324 13348 10885 13376
rect 8444 13336 8450 13348
rect 6730 13268 6736 13320
rect 6788 13308 6794 13320
rect 6917 13311 6975 13317
rect 6788 13280 6833 13308
rect 6788 13268 6794 13280
rect 6917 13277 6929 13311
rect 6963 13277 6975 13311
rect 6917 13271 6975 13277
rect 6932 13172 6960 13271
rect 7374 13268 7380 13320
rect 7432 13308 7438 13320
rect 8941 13311 8999 13317
rect 8941 13308 8953 13311
rect 7432 13280 8953 13308
rect 7432 13268 7438 13280
rect 8941 13277 8953 13280
rect 8987 13277 8999 13311
rect 9122 13308 9128 13320
rect 9083 13280 9128 13308
rect 8941 13271 8999 13277
rect 9122 13268 9128 13280
rect 9180 13268 9186 13320
rect 9232 13317 9260 13348
rect 10873 13345 10885 13348
rect 10919 13345 10931 13379
rect 10873 13339 10931 13345
rect 9217 13311 9275 13317
rect 9217 13277 9229 13311
rect 9263 13277 9275 13311
rect 9217 13271 9275 13277
rect 9309 13311 9367 13317
rect 9309 13277 9321 13311
rect 9355 13277 9367 13311
rect 9309 13271 9367 13277
rect 10965 13311 11023 13317
rect 10965 13277 10977 13311
rect 11011 13308 11023 13311
rect 11624 13308 11652 13416
rect 11698 13336 11704 13388
rect 11756 13376 11762 13388
rect 13449 13379 13507 13385
rect 13449 13376 13461 13379
rect 11756 13348 12756 13376
rect 11756 13336 11762 13348
rect 11011 13280 11652 13308
rect 11011 13277 11023 13280
rect 10965 13271 11023 13277
rect 7392 13240 7420 13268
rect 7561 13243 7619 13249
rect 7561 13240 7573 13243
rect 7392 13212 7573 13240
rect 7561 13209 7573 13212
rect 7607 13209 7619 13243
rect 7561 13203 7619 13209
rect 8297 13243 8355 13249
rect 8297 13209 8309 13243
rect 8343 13240 8355 13243
rect 8478 13240 8484 13252
rect 8343 13212 8484 13240
rect 8343 13209 8355 13212
rect 8297 13203 8355 13209
rect 8478 13200 8484 13212
rect 8536 13200 8542 13252
rect 8573 13243 8631 13249
rect 8573 13209 8585 13243
rect 8619 13240 8631 13243
rect 8754 13240 8760 13252
rect 8619 13212 8760 13240
rect 8619 13209 8631 13212
rect 8573 13203 8631 13209
rect 8754 13200 8760 13212
rect 8812 13200 8818 13252
rect 9324 13240 9352 13271
rect 12066 13268 12072 13320
rect 12124 13308 12130 13320
rect 12618 13317 12624 13320
rect 12437 13311 12495 13317
rect 12437 13308 12449 13311
rect 12124 13280 12449 13308
rect 12124 13268 12130 13280
rect 12437 13277 12449 13280
rect 12483 13277 12495 13311
rect 12437 13271 12495 13277
rect 12585 13311 12624 13317
rect 12585 13277 12597 13311
rect 12585 13271 12624 13277
rect 12618 13268 12624 13271
rect 12676 13268 12682 13320
rect 12728 13317 12756 13348
rect 13188 13348 13461 13376
rect 12713 13311 12771 13317
rect 12713 13277 12725 13311
rect 12759 13277 12771 13311
rect 12713 13271 12771 13277
rect 12943 13311 13001 13317
rect 12943 13277 12955 13311
rect 12989 13308 13001 13311
rect 13188 13308 13216 13348
rect 13449 13345 13461 13348
rect 13495 13345 13507 13379
rect 13740 13376 13768 13416
rect 13814 13404 13820 13456
rect 13872 13444 13878 13456
rect 14553 13447 14611 13453
rect 14553 13444 14565 13447
rect 13872 13416 14565 13444
rect 13872 13404 13878 13416
rect 14553 13413 14565 13416
rect 14599 13444 14611 13447
rect 14734 13444 14740 13456
rect 14599 13416 14740 13444
rect 14599 13413 14611 13416
rect 14553 13407 14611 13413
rect 14734 13404 14740 13416
rect 14792 13404 14798 13456
rect 16209 13447 16267 13453
rect 16209 13413 16221 13447
rect 16255 13444 16267 13447
rect 16666 13444 16672 13456
rect 16255 13416 16672 13444
rect 16255 13413 16267 13416
rect 16209 13407 16267 13413
rect 16666 13404 16672 13416
rect 16724 13404 16730 13456
rect 16022 13376 16028 13388
rect 13740 13348 16028 13376
rect 13449 13339 13507 13345
rect 16022 13336 16028 13348
rect 16080 13336 16086 13388
rect 16114 13336 16120 13388
rect 16172 13376 16178 13388
rect 16485 13379 16543 13385
rect 16485 13376 16497 13379
rect 16172 13348 16497 13376
rect 16172 13336 16178 13348
rect 16485 13345 16497 13348
rect 16531 13376 16543 13379
rect 16850 13376 16856 13388
rect 16531 13348 16856 13376
rect 16531 13345 16543 13348
rect 16485 13339 16543 13345
rect 16850 13336 16856 13348
rect 16908 13376 16914 13388
rect 17144 13376 17172 13484
rect 17954 13472 17960 13484
rect 18012 13472 18018 13524
rect 18693 13515 18751 13521
rect 18693 13481 18705 13515
rect 18739 13512 18751 13515
rect 20070 13512 20076 13524
rect 18739 13484 20076 13512
rect 18739 13481 18751 13484
rect 18693 13475 18751 13481
rect 20070 13472 20076 13484
rect 20128 13512 20134 13524
rect 20530 13512 20536 13524
rect 20128 13484 20536 13512
rect 20128 13472 20134 13484
rect 20530 13472 20536 13484
rect 20588 13472 20594 13524
rect 22002 13472 22008 13524
rect 22060 13512 22066 13524
rect 22189 13515 22247 13521
rect 22189 13512 22201 13515
rect 22060 13484 22201 13512
rect 22060 13472 22066 13484
rect 22189 13481 22201 13484
rect 22235 13481 22247 13515
rect 23842 13512 23848 13524
rect 23803 13484 23848 13512
rect 22189 13475 22247 13481
rect 23842 13472 23848 13484
rect 23900 13472 23906 13524
rect 24946 13472 24952 13524
rect 25004 13512 25010 13524
rect 25225 13515 25283 13521
rect 25225 13512 25237 13515
rect 25004 13484 25237 13512
rect 25004 13472 25010 13484
rect 25225 13481 25237 13484
rect 25271 13481 25283 13515
rect 25225 13475 25283 13481
rect 20898 13444 20904 13456
rect 16908 13348 17172 13376
rect 17236 13416 20904 13444
rect 16908 13336 16914 13348
rect 13354 13308 13360 13320
rect 12989 13280 13216 13308
rect 13315 13280 13360 13308
rect 12989 13277 13001 13280
rect 12943 13271 13001 13277
rect 13354 13268 13360 13280
rect 13412 13268 13418 13320
rect 13630 13268 13636 13320
rect 13688 13308 13694 13320
rect 14093 13311 14151 13317
rect 14093 13308 14105 13311
rect 13688 13280 14105 13308
rect 13688 13268 13694 13280
rect 14093 13277 14105 13280
rect 14139 13277 14151 13311
rect 14093 13271 14151 13277
rect 14277 13311 14335 13317
rect 14277 13277 14289 13311
rect 14323 13308 14335 13311
rect 15562 13308 15568 13320
rect 14323 13280 15568 13308
rect 14323 13277 14335 13280
rect 14277 13271 14335 13277
rect 15562 13268 15568 13280
rect 15620 13268 15626 13320
rect 15746 13308 15752 13320
rect 15707 13280 15752 13308
rect 15746 13268 15752 13280
rect 15804 13268 15810 13320
rect 16390 13308 16396 13320
rect 16351 13280 16396 13308
rect 16390 13268 16396 13280
rect 16448 13268 16454 13320
rect 16574 13268 16580 13320
rect 16632 13308 16638 13320
rect 17236 13317 17264 13416
rect 20898 13404 20904 13416
rect 20956 13404 20962 13456
rect 18046 13336 18052 13388
rect 18104 13376 18110 13388
rect 20993 13379 21051 13385
rect 20993 13376 21005 13379
rect 18104 13348 21005 13376
rect 18104 13336 18110 13348
rect 20993 13345 21005 13348
rect 21039 13345 21051 13379
rect 20993 13339 21051 13345
rect 22278 13336 22284 13388
rect 22336 13376 22342 13388
rect 22741 13379 22799 13385
rect 22741 13376 22753 13379
rect 22336 13348 22753 13376
rect 22336 13336 22342 13348
rect 22741 13345 22753 13348
rect 22787 13376 22799 13379
rect 23382 13376 23388 13388
rect 22787 13348 23388 13376
rect 22787 13345 22799 13348
rect 22741 13339 22799 13345
rect 23382 13336 23388 13348
rect 23440 13376 23446 13388
rect 24581 13379 24639 13385
rect 24581 13376 24593 13379
rect 23440 13348 24593 13376
rect 23440 13336 23446 13348
rect 24581 13345 24593 13348
rect 24627 13376 24639 13379
rect 24946 13376 24952 13388
rect 24627 13348 24952 13376
rect 24627 13345 24639 13348
rect 24581 13339 24639 13345
rect 24946 13336 24952 13348
rect 25004 13336 25010 13388
rect 16669 13311 16727 13317
rect 16669 13308 16681 13311
rect 16632 13280 16681 13308
rect 16632 13268 16638 13280
rect 16669 13277 16681 13280
rect 16715 13277 16727 13311
rect 16669 13271 16727 13277
rect 17221 13311 17279 13317
rect 17221 13277 17233 13311
rect 17267 13277 17279 13311
rect 17402 13308 17408 13320
rect 17363 13280 17408 13308
rect 17221 13271 17279 13277
rect 17402 13268 17408 13280
rect 17460 13268 17466 13320
rect 17497 13311 17555 13317
rect 17497 13277 17509 13311
rect 17543 13277 17555 13311
rect 17497 13271 17555 13277
rect 10226 13240 10232 13252
rect 9324 13212 10232 13240
rect 10226 13200 10232 13212
rect 10284 13200 10290 13252
rect 12805 13243 12863 13249
rect 12805 13209 12817 13243
rect 12851 13240 12863 13243
rect 14182 13240 14188 13252
rect 12851 13212 14188 13240
rect 12851 13209 12863 13212
rect 12805 13203 12863 13209
rect 14182 13200 14188 13212
rect 14240 13200 14246 13252
rect 17034 13240 17040 13252
rect 14292 13212 17040 13240
rect 7361 13175 7419 13181
rect 7361 13172 7373 13175
rect 6932 13144 7373 13172
rect 7361 13141 7373 13144
rect 7407 13172 7419 13175
rect 7466 13172 7472 13184
rect 7407 13144 7472 13172
rect 7407 13141 7419 13144
rect 7361 13135 7419 13141
rect 7466 13132 7472 13144
rect 7524 13132 7530 13184
rect 8202 13172 8208 13184
rect 8163 13144 8208 13172
rect 8202 13132 8208 13144
rect 8260 13132 8266 13184
rect 8389 13175 8447 13181
rect 8389 13141 8401 13175
rect 8435 13172 8447 13175
rect 8846 13172 8852 13184
rect 8435 13144 8852 13172
rect 8435 13141 8447 13144
rect 8389 13135 8447 13141
rect 8846 13132 8852 13144
rect 8904 13132 8910 13184
rect 8938 13132 8944 13184
rect 8996 13172 9002 13184
rect 9861 13175 9919 13181
rect 9861 13172 9873 13175
rect 8996 13144 9873 13172
rect 8996 13132 9002 13144
rect 9861 13141 9873 13144
rect 9907 13141 9919 13175
rect 9861 13135 9919 13141
rect 10029 13175 10087 13181
rect 10029 13141 10041 13175
rect 10075 13172 10087 13175
rect 11146 13172 11152 13184
rect 10075 13144 11152 13172
rect 10075 13141 10087 13144
rect 10029 13135 10087 13141
rect 11146 13132 11152 13144
rect 11204 13132 11210 13184
rect 12894 13132 12900 13184
rect 12952 13172 12958 13184
rect 13081 13175 13139 13181
rect 13081 13172 13093 13175
rect 12952 13144 13093 13172
rect 12952 13132 12958 13144
rect 13081 13141 13093 13144
rect 13127 13141 13139 13175
rect 13081 13135 13139 13141
rect 13170 13132 13176 13184
rect 13228 13172 13234 13184
rect 14292 13172 14320 13212
rect 17034 13200 17040 13212
rect 17092 13200 17098 13252
rect 15930 13172 15936 13184
rect 13228 13144 14320 13172
rect 15891 13144 15936 13172
rect 13228 13132 13234 13144
rect 15930 13132 15936 13144
rect 15988 13132 15994 13184
rect 17218 13132 17224 13184
rect 17276 13172 17282 13184
rect 17512 13172 17540 13271
rect 17586 13268 17592 13320
rect 17644 13308 17650 13320
rect 18233 13311 18291 13317
rect 17644 13280 17689 13308
rect 17644 13268 17650 13280
rect 18233 13277 18245 13311
rect 18279 13308 18291 13311
rect 18414 13308 18420 13320
rect 18279 13280 18420 13308
rect 18279 13277 18291 13280
rect 18233 13271 18291 13277
rect 18414 13268 18420 13280
rect 18472 13268 18478 13320
rect 18598 13308 18604 13320
rect 18559 13280 18604 13308
rect 18598 13268 18604 13280
rect 18656 13268 18662 13320
rect 18877 13311 18935 13317
rect 18877 13277 18889 13311
rect 18923 13308 18935 13311
rect 19242 13308 19248 13320
rect 18923 13280 19248 13308
rect 18923 13277 18935 13280
rect 18877 13271 18935 13277
rect 19242 13268 19248 13280
rect 19300 13268 19306 13320
rect 19521 13311 19579 13317
rect 19521 13277 19533 13311
rect 19567 13277 19579 13311
rect 19521 13271 19579 13277
rect 17954 13200 17960 13252
rect 18012 13240 18018 13252
rect 19536 13240 19564 13271
rect 19886 13268 19892 13320
rect 19944 13308 19950 13320
rect 20533 13311 20591 13317
rect 20533 13308 20545 13311
rect 19944 13280 20545 13308
rect 19944 13268 19950 13280
rect 20533 13277 20545 13280
rect 20579 13277 20591 13311
rect 21174 13308 21180 13320
rect 21135 13280 21180 13308
rect 20533 13271 20591 13277
rect 21174 13268 21180 13280
rect 21232 13268 21238 13320
rect 21545 13311 21603 13317
rect 21545 13277 21557 13311
rect 21591 13308 21603 13311
rect 21726 13308 21732 13320
rect 21591 13280 21732 13308
rect 21591 13277 21603 13280
rect 21545 13271 21603 13277
rect 21726 13268 21732 13280
rect 21784 13268 21790 13320
rect 22462 13268 22468 13320
rect 22520 13308 22526 13320
rect 22557 13311 22615 13317
rect 22557 13308 22569 13311
rect 22520 13280 22569 13308
rect 22520 13268 22526 13280
rect 22557 13277 22569 13280
rect 22603 13308 22615 13311
rect 23290 13308 23296 13320
rect 22603 13280 23296 13308
rect 22603 13277 22615 13280
rect 22557 13271 22615 13277
rect 23290 13268 23296 13280
rect 23348 13268 23354 13320
rect 23477 13311 23535 13317
rect 23477 13277 23489 13311
rect 23523 13277 23535 13311
rect 23658 13308 23664 13320
rect 23619 13280 23664 13308
rect 23477 13271 23535 13277
rect 20346 13240 20352 13252
rect 18012 13212 19564 13240
rect 20307 13212 20352 13240
rect 18012 13200 18018 13212
rect 20346 13200 20352 13212
rect 20404 13200 20410 13252
rect 23492 13240 23520 13271
rect 23658 13268 23664 13280
rect 23716 13268 23722 13320
rect 23934 13268 23940 13320
rect 23992 13308 23998 13320
rect 24762 13308 24768 13320
rect 23992 13280 24768 13308
rect 23992 13268 23998 13280
rect 24762 13268 24768 13280
rect 24820 13308 24826 13320
rect 25501 13311 25559 13317
rect 25501 13308 25513 13311
rect 24820 13280 25513 13308
rect 24820 13268 24826 13280
rect 25501 13277 25513 13280
rect 25547 13277 25559 13311
rect 25501 13271 25559 13277
rect 24670 13240 24676 13252
rect 20548 13212 21220 13240
rect 17276 13144 17540 13172
rect 17865 13175 17923 13181
rect 17276 13132 17282 13144
rect 17865 13141 17877 13175
rect 17911 13172 17923 13175
rect 18322 13172 18328 13184
rect 17911 13144 18328 13172
rect 17911 13141 17923 13144
rect 17865 13135 17923 13141
rect 18322 13132 18328 13144
rect 18380 13132 18386 13184
rect 18417 13175 18475 13181
rect 18417 13141 18429 13175
rect 18463 13172 18475 13175
rect 20548 13172 20576 13212
rect 21192 13184 21220 13212
rect 22066 13212 24676 13240
rect 20714 13172 20720 13184
rect 18463 13144 20576 13172
rect 20675 13144 20720 13172
rect 18463 13141 18475 13144
rect 18417 13135 18475 13141
rect 20714 13132 20720 13144
rect 20772 13132 20778 13184
rect 21174 13132 21180 13184
rect 21232 13132 21238 13184
rect 21634 13132 21640 13184
rect 21692 13172 21698 13184
rect 21729 13175 21787 13181
rect 21729 13172 21741 13175
rect 21692 13144 21741 13172
rect 21692 13132 21698 13144
rect 21729 13141 21741 13144
rect 21775 13172 21787 13175
rect 22066 13172 22094 13212
rect 24670 13200 24676 13212
rect 24728 13200 24734 13252
rect 24780 13212 25544 13240
rect 21775 13144 22094 13172
rect 21775 13141 21787 13144
rect 21729 13135 21787 13141
rect 22646 13132 22652 13184
rect 22704 13172 22710 13184
rect 24780 13181 24808 13212
rect 24765 13175 24823 13181
rect 22704 13144 22749 13172
rect 22704 13132 22710 13144
rect 24765 13141 24777 13175
rect 24811 13141 24823 13175
rect 24765 13135 24823 13141
rect 24854 13132 24860 13184
rect 24912 13172 24918 13184
rect 25314 13172 25320 13184
rect 24912 13144 25320 13172
rect 24912 13132 24918 13144
rect 25314 13132 25320 13144
rect 25372 13132 25378 13184
rect 25516 13172 25544 13212
rect 25590 13200 25596 13252
rect 25648 13240 25654 13252
rect 25746 13243 25804 13249
rect 25746 13240 25758 13243
rect 25648 13212 25758 13240
rect 25648 13200 25654 13212
rect 25746 13209 25758 13212
rect 25792 13209 25804 13243
rect 25746 13203 25804 13209
rect 25866 13172 25872 13184
rect 25516 13144 25872 13172
rect 25866 13132 25872 13144
rect 25924 13172 25930 13184
rect 26881 13175 26939 13181
rect 26881 13172 26893 13175
rect 25924 13144 26893 13172
rect 25924 13132 25930 13144
rect 26881 13141 26893 13144
rect 26927 13141 26939 13175
rect 26881 13135 26939 13141
rect 1104 13082 28888 13104
rect 1104 13030 10214 13082
rect 10266 13030 10278 13082
rect 10330 13030 10342 13082
rect 10394 13030 10406 13082
rect 10458 13030 10470 13082
rect 10522 13030 19478 13082
rect 19530 13030 19542 13082
rect 19594 13030 19606 13082
rect 19658 13030 19670 13082
rect 19722 13030 19734 13082
rect 19786 13030 28888 13082
rect 1104 13008 28888 13030
rect 6730 12928 6736 12980
rect 6788 12968 6794 12980
rect 6993 12971 7051 12977
rect 6993 12968 7005 12971
rect 6788 12940 7005 12968
rect 6788 12928 6794 12940
rect 6993 12937 7005 12940
rect 7039 12968 7051 12971
rect 7466 12968 7472 12980
rect 7039 12940 7328 12968
rect 7427 12940 7472 12968
rect 7039 12937 7051 12940
rect 6993 12931 7051 12937
rect 7098 12860 7104 12912
rect 7156 12900 7162 12912
rect 7193 12903 7251 12909
rect 7193 12900 7205 12903
rect 7156 12872 7205 12900
rect 7156 12860 7162 12872
rect 7193 12869 7205 12872
rect 7239 12869 7251 12903
rect 7300 12900 7328 12940
rect 7466 12928 7472 12940
rect 7524 12928 7530 12980
rect 7926 12968 7932 12980
rect 7887 12940 7932 12968
rect 7926 12928 7932 12940
rect 7984 12928 7990 12980
rect 8754 12928 8760 12980
rect 8812 12968 8818 12980
rect 9490 12968 9496 12980
rect 8812 12940 9496 12968
rect 8812 12928 8818 12940
rect 9490 12928 9496 12940
rect 9548 12928 9554 12980
rect 12526 12928 12532 12980
rect 12584 12968 12590 12980
rect 13173 12971 13231 12977
rect 13173 12968 13185 12971
rect 12584 12940 13185 12968
rect 12584 12928 12590 12940
rect 13173 12937 13185 12940
rect 13219 12968 13231 12971
rect 13630 12968 13636 12980
rect 13219 12940 13636 12968
rect 13219 12937 13231 12940
rect 13173 12931 13231 12937
rect 13630 12928 13636 12940
rect 13688 12928 13694 12980
rect 15654 12968 15660 12980
rect 15567 12940 15660 12968
rect 15654 12928 15660 12940
rect 15712 12968 15718 12980
rect 16942 12968 16948 12980
rect 15712 12940 16948 12968
rect 15712 12928 15718 12940
rect 16942 12928 16948 12940
rect 17000 12928 17006 12980
rect 17129 12971 17187 12977
rect 17129 12937 17141 12971
rect 17175 12968 17187 12971
rect 17402 12968 17408 12980
rect 17175 12940 17408 12968
rect 17175 12937 17187 12940
rect 17129 12931 17187 12937
rect 17402 12928 17408 12940
rect 17460 12928 17466 12980
rect 18325 12971 18383 12977
rect 18325 12937 18337 12971
rect 18371 12968 18383 12971
rect 18966 12968 18972 12980
rect 18371 12940 18972 12968
rect 18371 12937 18383 12940
rect 18325 12931 18383 12937
rect 18966 12928 18972 12940
rect 19024 12928 19030 12980
rect 19242 12928 19248 12980
rect 19300 12968 19306 12980
rect 19429 12971 19487 12977
rect 19429 12968 19441 12971
rect 19300 12940 19441 12968
rect 19300 12928 19306 12940
rect 19429 12937 19441 12940
rect 19475 12937 19487 12971
rect 19429 12931 19487 12937
rect 20438 12928 20444 12980
rect 20496 12968 20502 12980
rect 22738 12968 22744 12980
rect 20496 12940 22744 12968
rect 20496 12928 20502 12940
rect 22738 12928 22744 12940
rect 22796 12928 22802 12980
rect 24026 12968 24032 12980
rect 23987 12940 24032 12968
rect 24026 12928 24032 12940
rect 24084 12928 24090 12980
rect 25590 12968 25596 12980
rect 25551 12940 25596 12968
rect 25590 12928 25596 12940
rect 25648 12928 25654 12980
rect 8938 12909 8944 12912
rect 8909 12903 8944 12909
rect 8909 12900 8921 12903
rect 7300 12872 7696 12900
rect 7193 12863 7251 12869
rect 4430 12832 4436 12844
rect 4391 12804 4436 12832
rect 4430 12792 4436 12804
rect 4488 12792 4494 12844
rect 4700 12835 4758 12841
rect 4700 12801 4712 12835
rect 4746 12832 4758 12835
rect 5902 12832 5908 12844
rect 4746 12804 5908 12832
rect 4746 12801 4758 12804
rect 4700 12795 4758 12801
rect 5902 12792 5908 12804
rect 5960 12792 5966 12844
rect 7466 12832 7472 12844
rect 7427 12804 7472 12832
rect 7466 12792 7472 12804
rect 7524 12792 7530 12844
rect 7668 12841 7696 12872
rect 8128 12872 8921 12900
rect 8128 12841 8156 12872
rect 8909 12869 8921 12872
rect 8996 12900 9002 12912
rect 9125 12903 9183 12909
rect 8996 12872 9057 12900
rect 8909 12863 8944 12869
rect 8938 12860 8944 12863
rect 8996 12860 9002 12872
rect 9125 12869 9137 12903
rect 9171 12869 9183 12903
rect 12342 12900 12348 12912
rect 9125 12863 9183 12869
rect 11716 12872 12348 12900
rect 7653 12835 7711 12841
rect 7653 12801 7665 12835
rect 7699 12801 7711 12835
rect 7653 12795 7711 12801
rect 8113 12835 8171 12841
rect 8113 12801 8125 12835
rect 8159 12801 8171 12835
rect 8113 12795 8171 12801
rect 8297 12835 8355 12841
rect 8297 12801 8309 12835
rect 8343 12832 8355 12835
rect 8478 12832 8484 12844
rect 8343 12804 8484 12832
rect 8343 12801 8355 12804
rect 8297 12795 8355 12801
rect 7668 12696 7696 12795
rect 8478 12792 8484 12804
rect 8536 12792 8542 12844
rect 9140 12832 9168 12863
rect 11716 12841 11744 12872
rect 12342 12860 12348 12872
rect 12400 12900 12406 12912
rect 13725 12903 13783 12909
rect 13725 12900 13737 12903
rect 12400 12872 13737 12900
rect 12400 12860 12406 12872
rect 13725 12869 13737 12872
rect 13771 12869 13783 12903
rect 14366 12900 14372 12912
rect 14327 12872 14372 12900
rect 13725 12863 13783 12869
rect 14366 12860 14372 12872
rect 14424 12860 14430 12912
rect 15930 12900 15936 12912
rect 14844 12872 15936 12900
rect 11701 12835 11759 12841
rect 8680 12804 11468 12832
rect 8680 12776 8708 12804
rect 8018 12724 8024 12776
rect 8076 12764 8082 12776
rect 8205 12767 8263 12773
rect 8205 12764 8217 12767
rect 8076 12736 8217 12764
rect 8076 12724 8082 12736
rect 8205 12733 8217 12736
rect 8251 12733 8263 12767
rect 8205 12727 8263 12733
rect 8389 12767 8447 12773
rect 8389 12733 8401 12767
rect 8435 12764 8447 12767
rect 8662 12764 8668 12776
rect 8435 12736 8668 12764
rect 8435 12733 8447 12736
rect 8389 12727 8447 12733
rect 8662 12724 8668 12736
rect 8720 12724 8726 12776
rect 9674 12764 9680 12776
rect 8956 12736 9680 12764
rect 8757 12699 8815 12705
rect 8757 12696 8769 12699
rect 7668 12668 8769 12696
rect 8757 12665 8769 12668
rect 8803 12665 8815 12699
rect 8757 12659 8815 12665
rect 5813 12631 5871 12637
rect 5813 12597 5825 12631
rect 5859 12628 5871 12631
rect 6086 12628 6092 12640
rect 5859 12600 6092 12628
rect 5859 12597 5871 12600
rect 5813 12591 5871 12597
rect 6086 12588 6092 12600
rect 6144 12588 6150 12640
rect 6822 12628 6828 12640
rect 6783 12600 6828 12628
rect 6822 12588 6828 12600
rect 6880 12588 6886 12640
rect 7006 12628 7012 12640
rect 6967 12600 7012 12628
rect 7006 12588 7012 12600
rect 7064 12588 7070 12640
rect 8202 12588 8208 12640
rect 8260 12628 8266 12640
rect 8956 12637 8984 12736
rect 9674 12724 9680 12736
rect 9732 12724 9738 12776
rect 9858 12724 9864 12776
rect 9916 12764 9922 12776
rect 9953 12767 10011 12773
rect 9953 12764 9965 12767
rect 9916 12736 9965 12764
rect 9916 12724 9922 12736
rect 9953 12733 9965 12736
rect 9999 12733 10011 12767
rect 9953 12727 10011 12733
rect 11440 12696 11468 12804
rect 11701 12801 11713 12835
rect 11747 12801 11759 12835
rect 11701 12795 11759 12801
rect 12805 12835 12863 12841
rect 12805 12801 12817 12835
rect 12851 12832 12863 12835
rect 13170 12832 13176 12844
rect 12851 12804 13176 12832
rect 12851 12801 12863 12804
rect 12805 12795 12863 12801
rect 13170 12792 13176 12804
rect 13228 12792 13234 12844
rect 13265 12835 13323 12841
rect 13265 12801 13277 12835
rect 13311 12832 13323 12835
rect 14182 12832 14188 12844
rect 13311 12804 14188 12832
rect 13311 12801 13323 12804
rect 13265 12795 13323 12801
rect 14182 12792 14188 12804
rect 14240 12792 14246 12844
rect 14844 12841 14872 12872
rect 15930 12860 15936 12872
rect 15988 12900 15994 12912
rect 16390 12900 16396 12912
rect 15988 12872 16396 12900
rect 15988 12860 15994 12872
rect 16390 12860 16396 12872
rect 16448 12900 16454 12912
rect 16761 12903 16819 12909
rect 16761 12900 16773 12903
rect 16448 12872 16773 12900
rect 16448 12860 16454 12872
rect 16761 12869 16773 12872
rect 16807 12900 16819 12903
rect 16807 12872 17448 12900
rect 16807 12869 16819 12872
rect 16761 12863 16819 12869
rect 14553 12835 14611 12841
rect 14553 12801 14565 12835
rect 14599 12832 14611 12835
rect 14829 12835 14887 12841
rect 14829 12832 14841 12835
rect 14599 12804 14841 12832
rect 14599 12801 14611 12804
rect 14553 12795 14611 12801
rect 14829 12801 14841 12804
rect 14875 12801 14887 12835
rect 14829 12795 14887 12801
rect 15013 12835 15071 12841
rect 15013 12801 15025 12835
rect 15059 12801 15071 12835
rect 15013 12795 15071 12801
rect 11606 12764 11612 12776
rect 11567 12736 11612 12764
rect 11606 12724 11612 12736
rect 11664 12724 11670 12776
rect 12066 12764 12072 12776
rect 12027 12736 12072 12764
rect 12066 12724 12072 12736
rect 12124 12724 12130 12776
rect 13909 12767 13967 12773
rect 13909 12733 13921 12767
rect 13955 12764 13967 12767
rect 14458 12764 14464 12776
rect 13955 12736 14464 12764
rect 13955 12733 13967 12736
rect 13909 12727 13967 12733
rect 14458 12724 14464 12736
rect 14516 12764 14522 12776
rect 14642 12764 14648 12776
rect 14516 12736 14648 12764
rect 14516 12724 14522 12736
rect 14642 12724 14648 12736
rect 14700 12764 14706 12776
rect 15028 12764 15056 12795
rect 15286 12792 15292 12844
rect 15344 12832 15350 12844
rect 15838 12832 15844 12844
rect 15344 12804 15844 12832
rect 15344 12792 15350 12804
rect 15838 12792 15844 12804
rect 15896 12832 15902 12844
rect 16025 12835 16083 12841
rect 16025 12832 16037 12835
rect 15896 12804 16037 12832
rect 15896 12792 15902 12804
rect 16025 12801 16037 12804
rect 16071 12801 16083 12835
rect 16025 12795 16083 12801
rect 16117 12835 16175 12841
rect 16117 12801 16129 12835
rect 16163 12832 16175 12835
rect 16666 12832 16672 12844
rect 16163 12804 16672 12832
rect 16163 12801 16175 12804
rect 16117 12795 16175 12801
rect 16666 12792 16672 12804
rect 16724 12792 16730 12844
rect 17420 12841 17448 12872
rect 19168 12872 19840 12900
rect 16945 12835 17003 12841
rect 16945 12832 16957 12835
rect 16776 12804 16957 12832
rect 14700 12736 15056 12764
rect 15197 12767 15255 12773
rect 14700 12724 14706 12736
rect 15197 12733 15209 12767
rect 15243 12764 15255 12767
rect 15562 12764 15568 12776
rect 15243 12736 15568 12764
rect 15243 12733 15255 12736
rect 15197 12727 15255 12733
rect 15562 12724 15568 12736
rect 15620 12724 15626 12776
rect 13354 12696 13360 12708
rect 11440 12668 13360 12696
rect 13354 12656 13360 12668
rect 13412 12656 13418 12708
rect 14090 12656 14096 12708
rect 14148 12696 14154 12708
rect 16666 12696 16672 12708
rect 14148 12668 16672 12696
rect 14148 12656 14154 12668
rect 16666 12656 16672 12668
rect 16724 12696 16730 12708
rect 16776 12696 16804 12804
rect 16945 12801 16957 12804
rect 16991 12801 17003 12835
rect 16945 12795 17003 12801
rect 17405 12835 17463 12841
rect 17405 12801 17417 12835
rect 17451 12801 17463 12835
rect 17405 12795 17463 12801
rect 17494 12792 17500 12844
rect 17552 12832 17558 12844
rect 19168 12841 19196 12872
rect 19812 12841 19840 12872
rect 20898 12860 20904 12912
rect 20956 12900 20962 12912
rect 24578 12900 24584 12912
rect 20956 12872 24584 12900
rect 20956 12860 20962 12872
rect 24578 12860 24584 12872
rect 24636 12900 24642 12912
rect 24765 12903 24823 12909
rect 24765 12900 24777 12903
rect 24636 12872 24777 12900
rect 24636 12860 24642 12872
rect 24765 12869 24777 12872
rect 24811 12900 24823 12903
rect 26329 12903 26387 12909
rect 26329 12900 26341 12903
rect 24811 12872 26341 12900
rect 24811 12869 24823 12872
rect 24765 12863 24823 12869
rect 26329 12869 26341 12872
rect 26375 12869 26387 12903
rect 26329 12863 26387 12869
rect 17589 12835 17647 12841
rect 17589 12832 17601 12835
rect 17552 12804 17601 12832
rect 17552 12792 17558 12804
rect 17589 12801 17601 12804
rect 17635 12801 17647 12835
rect 17589 12795 17647 12801
rect 18233 12835 18291 12841
rect 18233 12801 18245 12835
rect 18279 12801 18291 12835
rect 18233 12795 18291 12801
rect 18417 12835 18475 12841
rect 18417 12801 18429 12835
rect 18463 12832 18475 12835
rect 19153 12835 19211 12841
rect 19153 12832 19165 12835
rect 18463 12804 19165 12832
rect 18463 12801 18475 12804
rect 18417 12795 18475 12801
rect 19153 12801 19165 12804
rect 19199 12801 19211 12835
rect 19153 12795 19211 12801
rect 19613 12835 19671 12841
rect 19613 12801 19625 12835
rect 19659 12801 19671 12835
rect 19613 12795 19671 12801
rect 19797 12835 19855 12841
rect 19797 12801 19809 12835
rect 19843 12832 19855 12835
rect 20162 12832 20168 12844
rect 19843 12804 20168 12832
rect 19843 12801 19855 12804
rect 19797 12795 19855 12801
rect 16850 12724 16856 12776
rect 16908 12764 16914 12776
rect 17512 12764 17540 12792
rect 16908 12736 17540 12764
rect 18248 12764 18276 12795
rect 18874 12764 18880 12776
rect 18248 12736 18880 12764
rect 16908 12724 16914 12736
rect 18874 12724 18880 12736
rect 18932 12724 18938 12776
rect 19334 12724 19340 12776
rect 19392 12724 19398 12776
rect 19352 12696 19380 12724
rect 16724 12668 16804 12696
rect 18708 12668 19380 12696
rect 16724 12656 16730 12668
rect 8941 12631 8999 12637
rect 8941 12628 8953 12631
rect 8260 12600 8953 12628
rect 8260 12588 8266 12600
rect 8941 12597 8953 12600
rect 8987 12597 8999 12631
rect 10962 12628 10968 12640
rect 10923 12600 10968 12628
rect 8941 12591 8999 12597
rect 10962 12588 10968 12600
rect 11020 12628 11026 12640
rect 12710 12628 12716 12640
rect 11020 12600 12716 12628
rect 11020 12588 11026 12600
rect 12710 12588 12716 12600
rect 12768 12588 12774 12640
rect 14185 12631 14243 12637
rect 14185 12597 14197 12631
rect 14231 12628 14243 12631
rect 14642 12628 14648 12640
rect 14231 12600 14648 12628
rect 14231 12597 14243 12600
rect 14185 12591 14243 12597
rect 14642 12588 14648 12600
rect 14700 12588 14706 12640
rect 16114 12588 16120 12640
rect 16172 12628 16178 12640
rect 16301 12631 16359 12637
rect 16301 12628 16313 12631
rect 16172 12600 16313 12628
rect 16172 12588 16178 12600
rect 16301 12597 16313 12600
rect 16347 12597 16359 12631
rect 16301 12591 16359 12597
rect 16574 12588 16580 12640
rect 16632 12628 16638 12640
rect 17218 12628 17224 12640
rect 16632 12600 17224 12628
rect 16632 12588 16638 12600
rect 17218 12588 17224 12600
rect 17276 12588 17282 12640
rect 17310 12588 17316 12640
rect 17368 12628 17374 12640
rect 18708 12637 18736 12668
rect 17773 12631 17831 12637
rect 17773 12628 17785 12631
rect 17368 12600 17785 12628
rect 17368 12588 17374 12600
rect 17773 12597 17785 12600
rect 17819 12597 17831 12631
rect 17773 12591 17831 12597
rect 18693 12631 18751 12637
rect 18693 12597 18705 12631
rect 18739 12597 18751 12631
rect 18874 12628 18880 12640
rect 18835 12600 18880 12628
rect 18693 12591 18751 12597
rect 18874 12588 18880 12600
rect 18932 12628 18938 12640
rect 19334 12628 19340 12640
rect 18932 12600 19340 12628
rect 18932 12588 18938 12600
rect 19334 12588 19340 12600
rect 19392 12628 19398 12640
rect 19628 12628 19656 12795
rect 20162 12792 20168 12804
rect 20220 12792 20226 12844
rect 20340 12835 20398 12841
rect 20340 12801 20352 12835
rect 20386 12832 20398 12835
rect 21082 12832 21088 12844
rect 20386 12804 21088 12832
rect 20386 12801 20398 12804
rect 20340 12795 20398 12801
rect 21082 12792 21088 12804
rect 21140 12792 21146 12844
rect 21174 12792 21180 12844
rect 21232 12832 21238 12844
rect 21913 12835 21971 12841
rect 21913 12832 21925 12835
rect 21232 12804 21925 12832
rect 21232 12792 21238 12804
rect 21913 12801 21925 12804
rect 21959 12801 21971 12835
rect 21913 12795 21971 12801
rect 22640 12835 22698 12841
rect 22640 12801 22652 12835
rect 22686 12832 22698 12835
rect 23014 12832 23020 12844
rect 22686 12804 23020 12832
rect 22686 12801 22698 12804
rect 22640 12795 22698 12801
rect 23014 12792 23020 12804
rect 23072 12792 23078 12844
rect 25406 12832 25412 12844
rect 25367 12804 25412 12832
rect 25406 12792 25412 12804
rect 25464 12792 25470 12844
rect 26050 12832 26056 12844
rect 26011 12804 26056 12832
rect 26050 12792 26056 12804
rect 26108 12792 26114 12844
rect 20070 12764 20076 12776
rect 20031 12736 20076 12764
rect 20070 12724 20076 12736
rect 20128 12724 20134 12776
rect 22373 12767 22431 12773
rect 22373 12733 22385 12767
rect 22419 12733 22431 12767
rect 24854 12764 24860 12776
rect 24815 12736 24860 12764
rect 22373 12727 22431 12733
rect 22097 12699 22155 12705
rect 22097 12665 22109 12699
rect 22143 12696 22155 12699
rect 22278 12696 22284 12708
rect 22143 12668 22284 12696
rect 22143 12665 22155 12668
rect 22097 12659 22155 12665
rect 22278 12656 22284 12668
rect 22336 12656 22342 12708
rect 21450 12628 21456 12640
rect 19392 12600 19656 12628
rect 21411 12600 21456 12628
rect 19392 12588 19398 12600
rect 21450 12588 21456 12600
rect 21508 12588 21514 12640
rect 22388 12628 22416 12727
rect 24854 12724 24860 12736
rect 24912 12724 24918 12776
rect 24946 12724 24952 12776
rect 25004 12764 25010 12776
rect 25004 12736 25049 12764
rect 25004 12724 25010 12736
rect 23474 12628 23480 12640
rect 22388 12600 23480 12628
rect 23474 12588 23480 12600
rect 23532 12588 23538 12640
rect 23750 12628 23756 12640
rect 23711 12600 23756 12628
rect 23750 12588 23756 12600
rect 23808 12588 23814 12640
rect 24397 12631 24455 12637
rect 24397 12597 24409 12631
rect 24443 12628 24455 12631
rect 24578 12628 24584 12640
rect 24443 12600 24584 12628
rect 24443 12597 24455 12600
rect 24397 12591 24455 12597
rect 24578 12588 24584 12600
rect 24636 12588 24642 12640
rect 25682 12588 25688 12640
rect 25740 12628 25746 12640
rect 25869 12631 25927 12637
rect 25869 12628 25881 12631
rect 25740 12600 25881 12628
rect 25740 12588 25746 12600
rect 25869 12597 25881 12600
rect 25915 12597 25927 12631
rect 28350 12628 28356 12640
rect 28311 12600 28356 12628
rect 25869 12591 25927 12597
rect 28350 12588 28356 12600
rect 28408 12588 28414 12640
rect 1104 12538 28888 12560
rect 1104 12486 5582 12538
rect 5634 12486 5646 12538
rect 5698 12486 5710 12538
rect 5762 12486 5774 12538
rect 5826 12486 5838 12538
rect 5890 12486 14846 12538
rect 14898 12486 14910 12538
rect 14962 12486 14974 12538
rect 15026 12486 15038 12538
rect 15090 12486 15102 12538
rect 15154 12486 24110 12538
rect 24162 12486 24174 12538
rect 24226 12486 24238 12538
rect 24290 12486 24302 12538
rect 24354 12486 24366 12538
rect 24418 12486 28888 12538
rect 1104 12464 28888 12486
rect 5537 12427 5595 12433
rect 5537 12393 5549 12427
rect 5583 12424 5595 12427
rect 5902 12424 5908 12436
rect 5583 12396 5908 12424
rect 5583 12393 5595 12396
rect 5537 12387 5595 12393
rect 5902 12384 5908 12396
rect 5960 12384 5966 12436
rect 6733 12427 6791 12433
rect 6733 12393 6745 12427
rect 6779 12424 6791 12427
rect 6914 12424 6920 12436
rect 6779 12396 6920 12424
rect 6779 12393 6791 12396
rect 6733 12387 6791 12393
rect 6914 12384 6920 12396
rect 6972 12384 6978 12436
rect 7006 12384 7012 12436
rect 7064 12424 7070 12436
rect 8386 12424 8392 12436
rect 7064 12396 8392 12424
rect 7064 12384 7070 12396
rect 8386 12384 8392 12396
rect 8444 12384 8450 12436
rect 8570 12424 8576 12436
rect 8483 12396 8576 12424
rect 8570 12384 8576 12396
rect 8628 12424 8634 12436
rect 9125 12427 9183 12433
rect 9125 12424 9137 12427
rect 8628 12396 9137 12424
rect 8628 12384 8634 12396
rect 9125 12393 9137 12396
rect 9171 12393 9183 12427
rect 9125 12387 9183 12393
rect 9674 12384 9680 12436
rect 9732 12424 9738 12436
rect 9953 12427 10011 12433
rect 9953 12424 9965 12427
rect 9732 12396 9965 12424
rect 9732 12384 9738 12396
rect 9953 12393 9965 12396
rect 9999 12393 10011 12427
rect 10594 12424 10600 12436
rect 9953 12387 10011 12393
rect 10336 12396 10600 12424
rect 6638 12316 6644 12368
rect 6696 12356 6702 12368
rect 7374 12356 7380 12368
rect 6696 12328 7380 12356
rect 6696 12316 6702 12328
rect 7374 12316 7380 12328
rect 7432 12356 7438 12368
rect 8018 12356 8024 12368
rect 7432 12328 8024 12356
rect 7432 12316 7438 12328
rect 8018 12316 8024 12328
rect 8076 12316 8082 12368
rect 8110 12316 8116 12368
rect 8168 12356 8174 12368
rect 9858 12356 9864 12368
rect 8168 12328 9864 12356
rect 8168 12316 8174 12328
rect 6822 12288 6828 12300
rect 5920 12260 6828 12288
rect 5920 12229 5948 12260
rect 6822 12248 6828 12260
rect 6880 12248 6886 12300
rect 5813 12223 5871 12229
rect 5813 12189 5825 12223
rect 5859 12189 5871 12223
rect 5813 12183 5871 12189
rect 5905 12223 5963 12229
rect 5905 12189 5917 12223
rect 5951 12189 5963 12223
rect 5905 12183 5963 12189
rect 5828 12152 5856 12183
rect 5994 12180 6000 12232
rect 6052 12220 6058 12232
rect 6181 12223 6239 12229
rect 6052 12192 6097 12220
rect 6052 12180 6058 12192
rect 6181 12189 6193 12223
rect 6227 12220 6239 12223
rect 6638 12220 6644 12232
rect 6227 12192 6644 12220
rect 6227 12189 6239 12192
rect 6181 12183 6239 12189
rect 6638 12180 6644 12192
rect 6696 12180 6702 12232
rect 7558 12180 7564 12232
rect 7616 12220 7622 12232
rect 8312 12229 8340 12328
rect 9858 12316 9864 12328
rect 9916 12316 9922 12368
rect 10042 12316 10048 12368
rect 10100 12356 10106 12368
rect 10336 12356 10364 12396
rect 10594 12384 10600 12396
rect 10652 12424 10658 12436
rect 11606 12424 11612 12436
rect 10652 12396 11612 12424
rect 10652 12384 10658 12396
rect 11606 12384 11612 12396
rect 11664 12384 11670 12436
rect 12342 12424 12348 12436
rect 12303 12396 12348 12424
rect 12342 12384 12348 12396
rect 12400 12384 12406 12436
rect 15378 12384 15384 12436
rect 15436 12424 15442 12436
rect 16574 12424 16580 12436
rect 15436 12396 16580 12424
rect 15436 12384 15442 12396
rect 16574 12384 16580 12396
rect 16632 12384 16638 12436
rect 20346 12384 20352 12436
rect 20404 12424 20410 12436
rect 20441 12427 20499 12433
rect 20441 12424 20453 12427
rect 20404 12396 20453 12424
rect 20404 12384 20410 12396
rect 20441 12393 20453 12396
rect 20487 12393 20499 12427
rect 20441 12387 20499 12393
rect 21818 12384 21824 12436
rect 21876 12424 21882 12436
rect 23477 12427 23535 12433
rect 23477 12424 23489 12427
rect 21876 12396 23489 12424
rect 21876 12384 21882 12396
rect 23477 12393 23489 12396
rect 23523 12424 23535 12427
rect 23934 12424 23940 12436
rect 23523 12396 23940 12424
rect 23523 12393 23535 12396
rect 23477 12387 23535 12393
rect 23934 12384 23940 12396
rect 23992 12384 23998 12436
rect 24765 12427 24823 12433
rect 24765 12393 24777 12427
rect 24811 12424 24823 12427
rect 26050 12424 26056 12436
rect 24811 12396 26056 12424
rect 24811 12393 24823 12396
rect 24765 12387 24823 12393
rect 26050 12384 26056 12396
rect 26108 12384 26114 12436
rect 10100 12328 10364 12356
rect 10100 12316 10106 12328
rect 8846 12248 8852 12300
rect 8904 12288 8910 12300
rect 10336 12297 10364 12328
rect 14550 12316 14556 12368
rect 14608 12356 14614 12368
rect 14826 12356 14832 12368
rect 14608 12328 14832 12356
rect 14608 12316 14614 12328
rect 14826 12316 14832 12328
rect 14884 12316 14890 12368
rect 15396 12356 15424 12384
rect 17586 12356 17592 12368
rect 14936 12328 15516 12356
rect 10321 12291 10379 12297
rect 8904 12260 10272 12288
rect 8904 12248 8910 12260
rect 7929 12223 7987 12229
rect 7929 12220 7941 12223
rect 7616 12192 7941 12220
rect 7616 12180 7622 12192
rect 7929 12189 7941 12192
rect 7975 12189 7987 12223
rect 7929 12183 7987 12189
rect 8297 12223 8355 12229
rect 8297 12189 8309 12223
rect 8343 12189 8355 12223
rect 8297 12183 8355 12189
rect 8573 12223 8631 12229
rect 8573 12189 8585 12223
rect 8619 12220 8631 12223
rect 8864 12220 8892 12248
rect 8619 12192 8892 12220
rect 8619 12189 8631 12192
rect 8573 12183 8631 12189
rect 9674 12180 9680 12232
rect 9732 12220 9738 12232
rect 10137 12223 10195 12229
rect 10137 12220 10149 12223
rect 9732 12192 10149 12220
rect 9732 12180 9738 12192
rect 10137 12189 10149 12192
rect 10183 12189 10195 12223
rect 10244 12220 10272 12260
rect 10321 12257 10333 12291
rect 10367 12257 10379 12291
rect 11974 12288 11980 12300
rect 11935 12260 11980 12288
rect 10321 12251 10379 12257
rect 11974 12248 11980 12260
rect 12032 12248 12038 12300
rect 14936 12288 14964 12328
rect 14568 12260 14964 12288
rect 11146 12220 11152 12232
rect 10244 12192 11152 12220
rect 10137 12183 10195 12189
rect 11146 12180 11152 12192
rect 11204 12180 11210 12232
rect 11992 12220 12020 12248
rect 13630 12220 13636 12232
rect 11992 12192 13636 12220
rect 13630 12180 13636 12192
rect 13688 12220 13694 12232
rect 13725 12223 13783 12229
rect 13725 12220 13737 12223
rect 13688 12192 13737 12220
rect 13688 12180 13694 12192
rect 13725 12189 13737 12192
rect 13771 12189 13783 12223
rect 13725 12183 13783 12189
rect 13814 12180 13820 12232
rect 13872 12220 13878 12232
rect 14568 12229 14596 12260
rect 15194 12248 15200 12300
rect 15252 12288 15258 12300
rect 15252 12260 15424 12288
rect 15252 12248 15258 12260
rect 14461 12223 14519 12229
rect 14461 12220 14473 12223
rect 13872 12192 14473 12220
rect 13872 12180 13878 12192
rect 14461 12189 14473 12192
rect 14507 12189 14519 12223
rect 14461 12183 14519 12189
rect 14553 12223 14611 12229
rect 14553 12189 14565 12223
rect 14599 12189 14611 12223
rect 14553 12183 14611 12189
rect 14642 12180 14648 12232
rect 14700 12220 14706 12232
rect 14700 12192 14745 12220
rect 14700 12180 14706 12192
rect 14826 12180 14832 12232
rect 14884 12220 14890 12232
rect 15396 12229 15424 12260
rect 15488 12229 15516 12328
rect 16040 12328 17592 12356
rect 15381 12223 15439 12229
rect 14884 12192 15332 12220
rect 14884 12180 14890 12192
rect 6086 12152 6092 12164
rect 5828 12124 6092 12152
rect 6086 12112 6092 12124
rect 6144 12152 6150 12164
rect 6546 12152 6552 12164
rect 6144 12124 6552 12152
rect 6144 12112 6150 12124
rect 6546 12112 6552 12124
rect 6604 12112 6610 12164
rect 6730 12112 6736 12164
rect 6788 12161 6794 12164
rect 6788 12155 6807 12161
rect 6795 12121 6807 12155
rect 7466 12152 7472 12164
rect 7379 12124 7472 12152
rect 6788 12115 6807 12121
rect 6788 12112 6794 12115
rect 7466 12112 7472 12124
rect 7524 12152 7530 12164
rect 8202 12152 8208 12164
rect 7524 12124 8208 12152
rect 7524 12112 7530 12124
rect 8202 12112 8208 12124
rect 8260 12152 8266 12164
rect 8481 12155 8539 12161
rect 8481 12152 8493 12155
rect 8260 12124 8493 12152
rect 8260 12112 8266 12124
rect 8481 12121 8493 12124
rect 8527 12121 8539 12155
rect 9093 12155 9151 12161
rect 9093 12152 9105 12155
rect 8481 12115 8539 12121
rect 8588 12124 9105 12152
rect 6917 12087 6975 12093
rect 6917 12053 6929 12087
rect 6963 12084 6975 12087
rect 7006 12084 7012 12096
rect 6963 12056 7012 12084
rect 6963 12053 6975 12056
rect 6917 12047 6975 12053
rect 7006 12044 7012 12056
rect 7064 12044 7070 12096
rect 7561 12087 7619 12093
rect 7561 12053 7573 12087
rect 7607 12084 7619 12087
rect 7742 12084 7748 12096
rect 7607 12056 7748 12084
rect 7607 12053 7619 12056
rect 7561 12047 7619 12053
rect 7742 12044 7748 12056
rect 7800 12044 7806 12096
rect 8018 12044 8024 12096
rect 8076 12084 8082 12096
rect 8588 12084 8616 12124
rect 9093 12121 9105 12124
rect 9139 12121 9151 12155
rect 9306 12152 9312 12164
rect 9267 12124 9312 12152
rect 9093 12115 9151 12121
rect 9306 12112 9312 12124
rect 9364 12112 9370 12164
rect 10870 12112 10876 12164
rect 10928 12152 10934 12164
rect 11710 12155 11768 12161
rect 11710 12152 11722 12155
rect 10928 12124 11722 12152
rect 10928 12112 10934 12124
rect 11710 12121 11722 12124
rect 11756 12121 11768 12155
rect 11710 12115 11768 12121
rect 13480 12155 13538 12161
rect 13480 12121 13492 12155
rect 13526 12152 13538 12155
rect 15105 12155 15163 12161
rect 15105 12152 15117 12155
rect 13526 12124 15117 12152
rect 13526 12121 13538 12124
rect 13480 12115 13538 12121
rect 15105 12121 15117 12124
rect 15151 12121 15163 12155
rect 15304 12152 15332 12192
rect 15381 12189 15393 12223
rect 15427 12189 15439 12223
rect 15381 12183 15439 12189
rect 15473 12223 15531 12229
rect 15473 12189 15485 12223
rect 15519 12189 15531 12223
rect 15473 12183 15531 12189
rect 15562 12180 15568 12232
rect 15620 12220 15626 12232
rect 16040 12229 16068 12328
rect 17586 12316 17592 12328
rect 17644 12316 17650 12368
rect 25038 12356 25044 12368
rect 24228 12328 25044 12356
rect 17034 12288 17040 12300
rect 16316 12260 17040 12288
rect 15749 12223 15807 12229
rect 15620 12192 15665 12220
rect 15620 12180 15626 12192
rect 15749 12189 15761 12223
rect 15795 12189 15807 12223
rect 15749 12183 15807 12189
rect 16025 12223 16083 12229
rect 16025 12189 16037 12223
rect 16071 12189 16083 12223
rect 16025 12183 16083 12189
rect 15764 12152 15792 12183
rect 16114 12180 16120 12232
rect 16172 12220 16178 12232
rect 16316 12229 16344 12260
rect 17034 12248 17040 12260
rect 17092 12248 17098 12300
rect 17218 12248 17224 12300
rect 17276 12288 17282 12300
rect 21085 12291 21143 12297
rect 17276 12260 17448 12288
rect 17276 12248 17282 12260
rect 16301 12223 16359 12229
rect 16172 12192 16217 12220
rect 16172 12180 16178 12192
rect 16301 12189 16313 12223
rect 16347 12189 16359 12223
rect 16301 12183 16359 12189
rect 16390 12180 16396 12232
rect 16448 12220 16454 12232
rect 17129 12223 17187 12229
rect 16448 12192 16493 12220
rect 16448 12180 16454 12192
rect 17129 12189 17141 12223
rect 17175 12189 17187 12223
rect 17310 12220 17316 12232
rect 17271 12192 17316 12220
rect 17129 12183 17187 12189
rect 17144 12152 17172 12183
rect 17310 12180 17316 12192
rect 17368 12180 17374 12232
rect 17420 12229 17448 12260
rect 21085 12257 21097 12291
rect 21131 12288 21143 12291
rect 21174 12288 21180 12300
rect 21131 12260 21180 12288
rect 21131 12257 21143 12260
rect 21085 12251 21143 12257
rect 21174 12248 21180 12260
rect 21232 12248 21238 12300
rect 22186 12288 22192 12300
rect 21468 12260 22192 12288
rect 17405 12223 17463 12229
rect 17405 12189 17417 12223
rect 17451 12189 17463 12223
rect 17405 12183 17463 12189
rect 17494 12180 17500 12232
rect 17552 12220 17558 12232
rect 19705 12223 19763 12229
rect 17552 12192 17597 12220
rect 17552 12180 17558 12192
rect 19705 12189 19717 12223
rect 19751 12220 19763 12223
rect 19978 12220 19984 12232
rect 19751 12192 19984 12220
rect 19751 12189 19763 12192
rect 19705 12183 19763 12189
rect 19978 12180 19984 12192
rect 20036 12180 20042 12232
rect 20806 12220 20812 12232
rect 20719 12192 20812 12220
rect 20806 12180 20812 12192
rect 20864 12220 20870 12232
rect 21358 12220 21364 12232
rect 20864 12192 21364 12220
rect 20864 12180 20870 12192
rect 21358 12180 21364 12192
rect 21416 12220 21422 12232
rect 21468 12220 21496 12260
rect 22186 12248 22192 12260
rect 22244 12248 22250 12300
rect 22278 12248 22284 12300
rect 22336 12288 22342 12300
rect 22741 12291 22799 12297
rect 22741 12288 22753 12291
rect 22336 12260 22753 12288
rect 22336 12248 22342 12260
rect 22741 12257 22753 12260
rect 22787 12257 22799 12291
rect 24228 12288 24256 12328
rect 25038 12316 25044 12328
rect 25096 12316 25102 12368
rect 22741 12251 22799 12257
rect 23308 12260 24256 12288
rect 24397 12291 24455 12297
rect 21634 12220 21640 12232
rect 21416 12192 21496 12220
rect 21595 12192 21640 12220
rect 21416 12180 21422 12192
rect 21634 12180 21640 12192
rect 21692 12180 21698 12232
rect 23308 12229 23336 12260
rect 24397 12257 24409 12291
rect 24443 12288 24455 12291
rect 24670 12288 24676 12300
rect 24443 12260 24676 12288
rect 24443 12257 24455 12260
rect 24397 12251 24455 12257
rect 24670 12248 24676 12260
rect 24728 12248 24734 12300
rect 21729 12223 21787 12229
rect 21729 12189 21741 12223
rect 21775 12220 21787 12223
rect 23293 12223 23351 12229
rect 21775 12192 22094 12220
rect 21775 12189 21787 12192
rect 21729 12183 21787 12189
rect 18046 12152 18052 12164
rect 15304 12124 18052 12152
rect 15105 12115 15163 12121
rect 18046 12112 18052 12124
rect 18104 12112 18110 12164
rect 19886 12152 19892 12164
rect 19847 12124 19892 12152
rect 19886 12112 19892 12124
rect 19944 12112 19950 12164
rect 8076 12056 8616 12084
rect 8076 12044 8082 12056
rect 8662 12044 8668 12096
rect 8720 12084 8726 12096
rect 8941 12087 8999 12093
rect 8941 12084 8953 12087
rect 8720 12056 8953 12084
rect 8720 12044 8726 12056
rect 8941 12053 8953 12056
rect 8987 12053 8999 12087
rect 14182 12084 14188 12096
rect 14143 12056 14188 12084
rect 8941 12047 8999 12053
rect 14182 12044 14188 12056
rect 14240 12044 14246 12096
rect 16574 12084 16580 12096
rect 16535 12056 16580 12084
rect 16574 12044 16580 12056
rect 16632 12044 16638 12096
rect 17770 12084 17776 12096
rect 17731 12056 17776 12084
rect 17770 12044 17776 12056
rect 17828 12044 17834 12096
rect 18233 12087 18291 12093
rect 18233 12053 18245 12087
rect 18279 12084 18291 12087
rect 18601 12087 18659 12093
rect 18601 12084 18613 12087
rect 18279 12056 18613 12084
rect 18279 12053 18291 12056
rect 18233 12047 18291 12053
rect 18601 12053 18613 12056
rect 18647 12084 18659 12087
rect 19334 12084 19340 12096
rect 18647 12056 19340 12084
rect 18647 12053 18659 12056
rect 18601 12047 18659 12053
rect 19334 12044 19340 12056
rect 19392 12044 19398 12096
rect 20901 12087 20959 12093
rect 20901 12053 20913 12087
rect 20947 12084 20959 12087
rect 21450 12084 21456 12096
rect 20947 12056 21456 12084
rect 20947 12053 20959 12056
rect 20901 12047 20959 12053
rect 21450 12044 21456 12056
rect 21508 12044 21514 12096
rect 21910 12084 21916 12096
rect 21871 12056 21916 12084
rect 21910 12044 21916 12056
rect 21968 12044 21974 12096
rect 22066 12084 22094 12192
rect 23293 12189 23305 12223
rect 23339 12189 23351 12223
rect 23293 12183 23351 12189
rect 23566 12180 23572 12232
rect 23624 12220 23630 12232
rect 23750 12220 23756 12232
rect 23624 12192 23756 12220
rect 23624 12180 23630 12192
rect 23750 12180 23756 12192
rect 23808 12180 23814 12232
rect 24026 12220 24032 12232
rect 23987 12192 24032 12220
rect 24026 12180 24032 12192
rect 24084 12180 24090 12232
rect 24578 12220 24584 12232
rect 24539 12192 24584 12220
rect 24578 12180 24584 12192
rect 24636 12180 24642 12232
rect 24762 12180 24768 12232
rect 24820 12220 24826 12232
rect 25409 12223 25467 12229
rect 25409 12220 25421 12223
rect 24820 12192 25421 12220
rect 24820 12180 24826 12192
rect 25409 12189 25421 12192
rect 25455 12220 25467 12223
rect 25455 12192 25544 12220
rect 25455 12189 25467 12192
rect 25409 12183 25467 12189
rect 22554 12152 22560 12164
rect 22467 12124 22560 12152
rect 22554 12112 22560 12124
rect 22612 12152 22618 12164
rect 25041 12155 25099 12161
rect 25041 12152 25053 12155
rect 22612 12124 25053 12152
rect 22612 12112 22618 12124
rect 25041 12121 25053 12124
rect 25087 12121 25099 12155
rect 25041 12115 25099 12121
rect 22189 12087 22247 12093
rect 22189 12084 22201 12087
rect 22066 12056 22201 12084
rect 22189 12053 22201 12056
rect 22235 12053 22247 12087
rect 22189 12047 22247 12053
rect 22649 12087 22707 12093
rect 22649 12053 22661 12087
rect 22695 12084 22707 12087
rect 23566 12084 23572 12096
rect 22695 12056 23572 12084
rect 22695 12053 22707 12056
rect 22649 12047 22707 12053
rect 23566 12044 23572 12056
rect 23624 12044 23630 12096
rect 23842 12084 23848 12096
rect 23803 12056 23848 12084
rect 23842 12044 23848 12056
rect 23900 12044 23906 12096
rect 25516 12084 25544 12192
rect 25682 12161 25688 12164
rect 25676 12115 25688 12161
rect 25740 12152 25746 12164
rect 25740 12124 25776 12152
rect 25682 12112 25688 12115
rect 25740 12112 25746 12124
rect 25774 12084 25780 12096
rect 25516 12056 25780 12084
rect 25774 12044 25780 12056
rect 25832 12044 25838 12096
rect 25958 12044 25964 12096
rect 26016 12084 26022 12096
rect 26789 12087 26847 12093
rect 26789 12084 26801 12087
rect 26016 12056 26801 12084
rect 26016 12044 26022 12056
rect 26789 12053 26801 12056
rect 26835 12053 26847 12087
rect 26789 12047 26847 12053
rect 1104 11994 28888 12016
rect 1104 11942 10214 11994
rect 10266 11942 10278 11994
rect 10330 11942 10342 11994
rect 10394 11942 10406 11994
rect 10458 11942 10470 11994
rect 10522 11942 19478 11994
rect 19530 11942 19542 11994
rect 19594 11942 19606 11994
rect 19658 11942 19670 11994
rect 19722 11942 19734 11994
rect 19786 11942 28888 11994
rect 1104 11920 28888 11942
rect 7098 11880 7104 11892
rect 5184 11852 7104 11880
rect 4522 11704 4528 11756
rect 4580 11744 4586 11756
rect 5184 11744 5212 11852
rect 6932 11821 6960 11852
rect 7098 11840 7104 11852
rect 7156 11840 7162 11892
rect 7834 11840 7840 11892
rect 7892 11880 7898 11892
rect 10686 11880 10692 11892
rect 7892 11852 10692 11880
rect 7892 11840 7898 11852
rect 10686 11840 10692 11852
rect 10744 11840 10750 11892
rect 10870 11880 10876 11892
rect 10831 11852 10876 11880
rect 10870 11840 10876 11852
rect 10928 11840 10934 11892
rect 11146 11840 11152 11892
rect 11204 11880 11210 11892
rect 12250 11880 12256 11892
rect 11204 11852 12256 11880
rect 11204 11840 11210 11852
rect 12250 11840 12256 11852
rect 12308 11840 12314 11892
rect 12986 11880 12992 11892
rect 12947 11852 12992 11880
rect 12986 11840 12992 11852
rect 13044 11840 13050 11892
rect 15838 11880 15844 11892
rect 15799 11852 15844 11880
rect 15838 11840 15844 11852
rect 15896 11840 15902 11892
rect 17862 11840 17868 11892
rect 17920 11880 17926 11892
rect 18325 11883 18383 11889
rect 18325 11880 18337 11883
rect 17920 11852 18337 11880
rect 17920 11840 17926 11852
rect 18325 11849 18337 11852
rect 18371 11849 18383 11883
rect 20438 11880 20444 11892
rect 18325 11843 18383 11849
rect 19306 11852 20444 11880
rect 5261 11815 5319 11821
rect 5261 11781 5273 11815
rect 5307 11812 5319 11815
rect 5813 11815 5871 11821
rect 5813 11812 5825 11815
rect 5307 11784 5825 11812
rect 5307 11781 5319 11784
rect 5261 11775 5319 11781
rect 5813 11781 5825 11784
rect 5859 11781 5871 11815
rect 5813 11775 5871 11781
rect 6917 11815 6975 11821
rect 6917 11781 6929 11815
rect 6963 11781 6975 11815
rect 7466 11812 7472 11824
rect 6917 11775 6975 11781
rect 7024 11784 7472 11812
rect 5353 11747 5411 11753
rect 5353 11744 5365 11747
rect 4580 11716 5365 11744
rect 4580 11704 4586 11716
rect 5353 11713 5365 11716
rect 5399 11713 5411 11747
rect 5353 11707 5411 11713
rect 5629 11747 5687 11753
rect 5629 11713 5641 11747
rect 5675 11713 5687 11747
rect 5629 11707 5687 11713
rect 5905 11747 5963 11753
rect 5905 11713 5917 11747
rect 5951 11744 5963 11747
rect 5994 11744 6000 11756
rect 5951 11716 6000 11744
rect 5951 11713 5963 11716
rect 5905 11707 5963 11713
rect 5644 11676 5672 11707
rect 5994 11704 6000 11716
rect 6052 11744 6058 11756
rect 6733 11747 6791 11753
rect 6052 11716 6684 11744
rect 6052 11704 6058 11716
rect 5644 11648 6592 11676
rect 6564 11617 6592 11648
rect 6549 11611 6607 11617
rect 6549 11577 6561 11611
rect 6595 11577 6607 11611
rect 6656 11608 6684 11716
rect 6733 11713 6745 11747
rect 6779 11713 6791 11747
rect 6733 11707 6791 11713
rect 6825 11747 6883 11753
rect 6825 11713 6837 11747
rect 6871 11744 6883 11747
rect 7024 11744 7052 11784
rect 7466 11772 7472 11784
rect 7524 11772 7530 11824
rect 14182 11772 14188 11824
rect 14240 11812 14246 11824
rect 14338 11815 14396 11821
rect 14338 11812 14350 11815
rect 14240 11784 14350 11812
rect 14240 11772 14246 11784
rect 14338 11781 14350 11784
rect 14384 11781 14396 11815
rect 15856 11812 15884 11840
rect 14338 11775 14396 11781
rect 14476 11784 15884 11812
rect 6871 11716 7052 11744
rect 7101 11747 7159 11753
rect 6871 11713 6883 11716
rect 6825 11707 6883 11713
rect 7101 11713 7113 11747
rect 7147 11713 7159 11747
rect 7101 11707 7159 11713
rect 7193 11747 7251 11753
rect 7193 11713 7205 11747
rect 7239 11744 7251 11747
rect 7374 11744 7380 11756
rect 7239 11716 7380 11744
rect 7239 11713 7251 11716
rect 7193 11707 7251 11713
rect 6748 11676 6776 11707
rect 7006 11676 7012 11688
rect 6748 11648 7012 11676
rect 7006 11636 7012 11648
rect 7064 11636 7070 11688
rect 7116 11676 7144 11707
rect 7374 11704 7380 11716
rect 7432 11744 7438 11756
rect 7650 11744 7656 11756
rect 7432 11716 7656 11744
rect 7432 11704 7438 11716
rect 7650 11704 7656 11716
rect 7708 11704 7714 11756
rect 7745 11747 7803 11753
rect 7745 11713 7757 11747
rect 7791 11744 7803 11747
rect 8386 11744 8392 11756
rect 7791 11716 8392 11744
rect 7791 11713 7803 11716
rect 7745 11707 7803 11713
rect 8386 11704 8392 11716
rect 8444 11704 8450 11756
rect 9309 11747 9367 11753
rect 9309 11713 9321 11747
rect 9355 11713 9367 11747
rect 9309 11707 9367 11713
rect 7558 11676 7564 11688
rect 7116 11648 7564 11676
rect 7558 11636 7564 11648
rect 7616 11636 7622 11688
rect 8021 11679 8079 11685
rect 8021 11645 8033 11679
rect 8067 11676 8079 11679
rect 8202 11676 8208 11688
rect 8067 11648 8208 11676
rect 8067 11645 8079 11648
rect 8021 11639 8079 11645
rect 8202 11636 8208 11648
rect 8260 11636 8266 11688
rect 8754 11636 8760 11688
rect 8812 11676 8818 11688
rect 9217 11679 9275 11685
rect 9217 11676 9229 11679
rect 8812 11648 9229 11676
rect 8812 11636 8818 11648
rect 9217 11645 9229 11648
rect 9263 11645 9275 11679
rect 9217 11639 9275 11645
rect 7650 11608 7656 11620
rect 6656 11580 7656 11608
rect 6549 11571 6607 11577
rect 7650 11568 7656 11580
rect 7708 11568 7714 11620
rect 9324 11608 9352 11707
rect 9674 11704 9680 11756
rect 9732 11744 9738 11756
rect 9769 11747 9827 11753
rect 9769 11744 9781 11747
rect 9732 11716 9781 11744
rect 9732 11704 9738 11716
rect 9769 11713 9781 11716
rect 9815 11713 9827 11747
rect 9769 11707 9827 11713
rect 9953 11747 10011 11753
rect 9953 11713 9965 11747
rect 9999 11744 10011 11747
rect 10042 11744 10048 11756
rect 9999 11716 10048 11744
rect 9999 11713 10011 11716
rect 9953 11707 10011 11713
rect 10042 11704 10048 11716
rect 10100 11704 10106 11756
rect 10226 11744 10232 11756
rect 10187 11716 10232 11744
rect 10226 11704 10232 11716
rect 10284 11704 10290 11756
rect 10318 11704 10324 11756
rect 10376 11728 10382 11756
rect 10413 11747 10471 11753
rect 10413 11728 10425 11747
rect 10376 11713 10425 11728
rect 10459 11713 10471 11747
rect 10376 11707 10471 11713
rect 10508 11750 10566 11756
rect 10508 11716 10520 11750
rect 10554 11716 10566 11750
rect 10508 11710 10566 11716
rect 10376 11704 10456 11707
rect 10336 11700 10456 11704
rect 10318 11608 10324 11620
rect 9324 11580 10324 11608
rect 10318 11568 10324 11580
rect 10376 11568 10382 11620
rect 5442 11500 5448 11552
rect 5500 11540 5506 11552
rect 5629 11543 5687 11549
rect 5629 11540 5641 11543
rect 5500 11512 5641 11540
rect 5500 11500 5506 11512
rect 5629 11509 5641 11512
rect 5675 11509 5687 11543
rect 5629 11503 5687 11509
rect 6822 11500 6828 11552
rect 6880 11540 6886 11552
rect 8941 11543 8999 11549
rect 8941 11540 8953 11543
rect 6880 11512 8953 11540
rect 6880 11500 6886 11512
rect 8941 11509 8953 11512
rect 8987 11509 8999 11543
rect 9766 11540 9772 11552
rect 9727 11512 9772 11540
rect 8941 11503 8999 11509
rect 9766 11500 9772 11512
rect 9824 11500 9830 11552
rect 10134 11500 10140 11552
rect 10192 11540 10198 11552
rect 10520 11540 10548 11710
rect 10594 11704 10600 11756
rect 10652 11744 10658 11756
rect 12066 11744 12072 11756
rect 10652 11716 10697 11744
rect 12027 11716 12072 11744
rect 10652 11704 10658 11716
rect 12066 11704 12072 11716
rect 12124 11704 12130 11756
rect 12250 11704 12256 11756
rect 12308 11744 12314 11756
rect 12529 11747 12587 11753
rect 12529 11744 12541 11747
rect 12308 11716 12541 11744
rect 12308 11704 12314 11716
rect 12529 11713 12541 11716
rect 12575 11713 12587 11747
rect 12529 11707 12587 11713
rect 12713 11747 12771 11753
rect 12713 11713 12725 11747
rect 12759 11713 12771 11747
rect 12713 11707 12771 11713
rect 12728 11676 12756 11707
rect 13630 11704 13636 11756
rect 13688 11744 13694 11756
rect 14093 11747 14151 11753
rect 14093 11744 14105 11747
rect 13688 11716 14105 11744
rect 13688 11704 13694 11716
rect 14093 11713 14105 11716
rect 14139 11713 14151 11747
rect 14476 11744 14504 11784
rect 16574 11772 16580 11824
rect 16632 11812 16638 11824
rect 17782 11815 17840 11821
rect 17782 11812 17794 11815
rect 16632 11784 17794 11812
rect 16632 11772 16638 11784
rect 17782 11781 17794 11784
rect 17828 11781 17840 11815
rect 19306 11812 19334 11852
rect 20438 11840 20444 11852
rect 20496 11880 20502 11892
rect 20898 11880 20904 11892
rect 20496 11852 20904 11880
rect 20496 11840 20502 11852
rect 20898 11840 20904 11852
rect 20956 11840 20962 11892
rect 21082 11880 21088 11892
rect 21043 11852 21088 11880
rect 21082 11840 21088 11852
rect 21140 11840 21146 11892
rect 23014 11880 23020 11892
rect 22066 11852 22876 11880
rect 22975 11852 23020 11880
rect 17782 11775 17840 11781
rect 18708 11784 19334 11812
rect 20533 11815 20591 11821
rect 14093 11707 14151 11713
rect 14200 11716 14504 11744
rect 13722 11676 13728 11688
rect 12728 11648 13728 11676
rect 13722 11636 13728 11648
rect 13780 11676 13786 11688
rect 14200 11676 14228 11716
rect 15286 11704 15292 11756
rect 15344 11744 15350 11756
rect 15933 11747 15991 11753
rect 15933 11744 15945 11747
rect 15344 11716 15945 11744
rect 15344 11704 15350 11716
rect 15933 11713 15945 11716
rect 15979 11713 15991 11747
rect 15933 11707 15991 11713
rect 13780 11648 14228 11676
rect 13780 11636 13786 11648
rect 11609 11611 11667 11617
rect 11609 11577 11621 11611
rect 11655 11608 11667 11611
rect 13170 11608 13176 11620
rect 11655 11580 13176 11608
rect 11655 11577 11667 11580
rect 11609 11571 11667 11577
rect 10192 11512 10548 11540
rect 10192 11500 10198 11512
rect 10594 11500 10600 11552
rect 10652 11540 10658 11552
rect 11624 11540 11652 11571
rect 13170 11568 13176 11580
rect 13228 11568 13234 11620
rect 15948 11608 15976 11707
rect 17034 11704 17040 11756
rect 17092 11744 17098 11756
rect 18708 11744 18736 11784
rect 20533 11781 20545 11815
rect 20579 11812 20591 11815
rect 20990 11812 20996 11824
rect 20579 11784 20996 11812
rect 20579 11781 20591 11784
rect 20533 11775 20591 11781
rect 20990 11772 20996 11784
rect 21048 11772 21054 11824
rect 21910 11772 21916 11824
rect 21968 11812 21974 11824
rect 22066 11812 22094 11852
rect 21968 11784 22094 11812
rect 21968 11772 21974 11784
rect 17092 11716 18736 11744
rect 18785 11747 18843 11753
rect 17092 11704 17098 11716
rect 18785 11713 18797 11747
rect 18831 11713 18843 11747
rect 18785 11707 18843 11713
rect 19521 11747 19579 11753
rect 19521 11713 19533 11747
rect 19567 11744 19579 11747
rect 19978 11744 19984 11756
rect 19567 11716 19984 11744
rect 19567 11713 19579 11716
rect 19521 11707 19579 11713
rect 18046 11676 18052 11688
rect 18007 11648 18052 11676
rect 18046 11636 18052 11648
rect 18104 11636 18110 11688
rect 18800 11676 18828 11707
rect 19978 11704 19984 11716
rect 20036 11704 20042 11756
rect 20714 11704 20720 11756
rect 20772 11744 20778 11756
rect 21269 11747 21327 11753
rect 21269 11744 21281 11747
rect 20772 11716 21281 11744
rect 20772 11704 20778 11716
rect 21269 11713 21281 11716
rect 21315 11713 21327 11747
rect 21269 11707 21327 11713
rect 22094 11704 22100 11756
rect 22152 11744 22158 11756
rect 22152 11716 22197 11744
rect 22152 11704 22158 11716
rect 22370 11704 22376 11756
rect 22428 11744 22434 11756
rect 22741 11747 22799 11753
rect 22741 11744 22753 11747
rect 22428 11716 22753 11744
rect 22428 11704 22434 11716
rect 22741 11713 22753 11716
rect 22787 11713 22799 11747
rect 22848 11744 22876 11852
rect 23014 11840 23020 11852
rect 23072 11840 23078 11892
rect 24486 11880 24492 11892
rect 24447 11852 24492 11880
rect 24486 11840 24492 11852
rect 24544 11840 24550 11892
rect 24854 11840 24860 11892
rect 24912 11880 24918 11892
rect 25958 11880 25964 11892
rect 24912 11852 25964 11880
rect 24912 11840 24918 11852
rect 25958 11840 25964 11852
rect 26016 11840 26022 11892
rect 23569 11815 23627 11821
rect 23569 11812 23581 11815
rect 23308 11784 23581 11812
rect 23201 11747 23259 11753
rect 23201 11744 23213 11747
rect 22848 11716 23213 11744
rect 22741 11707 22799 11713
rect 23201 11713 23213 11716
rect 23247 11713 23259 11747
rect 23201 11707 23259 11713
rect 20254 11676 20260 11688
rect 18800 11648 20260 11676
rect 20254 11636 20260 11648
rect 20312 11636 20318 11688
rect 20625 11679 20683 11685
rect 20625 11645 20637 11679
rect 20671 11676 20683 11679
rect 21174 11676 21180 11688
rect 20671 11648 21180 11676
rect 20671 11645 20683 11648
rect 20625 11639 20683 11645
rect 16669 11611 16727 11617
rect 16669 11608 16681 11611
rect 15948 11580 16681 11608
rect 16669 11577 16681 11580
rect 16715 11577 16727 11611
rect 16669 11571 16727 11577
rect 20530 11568 20536 11620
rect 20588 11608 20594 11620
rect 20640 11608 20668 11639
rect 21174 11636 21180 11648
rect 21232 11636 21238 11688
rect 22281 11679 22339 11685
rect 22281 11676 22293 11679
rect 22066 11648 22293 11676
rect 20588 11580 20668 11608
rect 20588 11568 20594 11580
rect 10652 11512 11652 11540
rect 10652 11500 10658 11512
rect 11974 11500 11980 11552
rect 12032 11540 12038 11552
rect 12161 11543 12219 11549
rect 12161 11540 12173 11543
rect 12032 11512 12173 11540
rect 12032 11500 12038 11512
rect 12161 11509 12173 11512
rect 12207 11509 12219 11543
rect 12161 11503 12219 11509
rect 12621 11543 12679 11549
rect 12621 11509 12633 11543
rect 12667 11540 12679 11543
rect 13262 11540 13268 11552
rect 12667 11512 13268 11540
rect 12667 11509 12679 11512
rect 12621 11503 12679 11509
rect 13262 11500 13268 11512
rect 13320 11500 13326 11552
rect 13814 11540 13820 11552
rect 13775 11512 13820 11540
rect 13814 11500 13820 11512
rect 13872 11500 13878 11552
rect 13906 11500 13912 11552
rect 13964 11540 13970 11552
rect 15473 11543 15531 11549
rect 15473 11540 15485 11543
rect 13964 11512 15485 11540
rect 13964 11500 13970 11512
rect 15473 11509 15485 11512
rect 15519 11509 15531 11543
rect 15473 11503 15531 11509
rect 16114 11500 16120 11552
rect 16172 11540 16178 11552
rect 18506 11540 18512 11552
rect 16172 11512 18512 11540
rect 16172 11500 16178 11512
rect 18506 11500 18512 11512
rect 18564 11500 18570 11552
rect 18966 11540 18972 11552
rect 18927 11512 18972 11540
rect 18966 11500 18972 11512
rect 19024 11500 19030 11552
rect 19150 11500 19156 11552
rect 19208 11540 19214 11552
rect 19337 11543 19395 11549
rect 19337 11540 19349 11543
rect 19208 11512 19349 11540
rect 19208 11500 19214 11512
rect 19337 11509 19349 11512
rect 19383 11509 19395 11543
rect 19337 11503 19395 11509
rect 20073 11543 20131 11549
rect 20073 11509 20085 11543
rect 20119 11540 20131 11543
rect 20346 11540 20352 11552
rect 20119 11512 20352 11540
rect 20119 11509 20131 11512
rect 20073 11503 20131 11509
rect 20346 11500 20352 11512
rect 20404 11500 20410 11552
rect 21174 11500 21180 11552
rect 21232 11540 21238 11552
rect 22066 11540 22094 11648
rect 22281 11645 22293 11648
rect 22327 11676 22339 11679
rect 23308 11676 23336 11784
rect 23569 11781 23581 11784
rect 23615 11781 23627 11815
rect 23569 11775 23627 11781
rect 23753 11815 23811 11821
rect 23753 11781 23765 11815
rect 23799 11812 23811 11815
rect 24762 11812 24768 11824
rect 23799 11784 24768 11812
rect 23799 11781 23811 11784
rect 23753 11775 23811 11781
rect 23474 11704 23480 11756
rect 23532 11744 23538 11756
rect 23768 11744 23796 11775
rect 24762 11772 24768 11784
rect 24820 11772 24826 11824
rect 25314 11772 25320 11824
rect 25372 11812 25378 11824
rect 28077 11815 28135 11821
rect 28077 11812 28089 11815
rect 25372 11784 28089 11812
rect 25372 11772 25378 11784
rect 28077 11781 28089 11784
rect 28123 11781 28135 11815
rect 28077 11775 28135 11781
rect 23532 11716 23796 11744
rect 24581 11747 24639 11753
rect 23532 11704 23538 11716
rect 24581 11713 24593 11747
rect 24627 11744 24639 11747
rect 25130 11744 25136 11756
rect 24627 11716 25136 11744
rect 24627 11713 24639 11716
rect 24581 11707 24639 11713
rect 25130 11704 25136 11716
rect 25188 11704 25194 11756
rect 27801 11747 27859 11753
rect 25516 11716 26188 11744
rect 25516 11688 25544 11716
rect 22327 11648 23336 11676
rect 24765 11679 24823 11685
rect 22327 11645 22339 11648
rect 22281 11639 22339 11645
rect 24765 11645 24777 11679
rect 24811 11676 24823 11679
rect 25498 11676 25504 11688
rect 24811 11648 25504 11676
rect 24811 11645 24823 11648
rect 24765 11639 24823 11645
rect 25498 11636 25504 11648
rect 25556 11636 25562 11688
rect 26050 11676 26056 11688
rect 26011 11648 26056 11676
rect 26050 11636 26056 11648
rect 26108 11636 26114 11688
rect 26160 11685 26188 11716
rect 27801 11713 27813 11747
rect 27847 11744 27859 11747
rect 28258 11744 28264 11756
rect 27847 11716 28264 11744
rect 27847 11713 27859 11716
rect 27801 11707 27859 11713
rect 28258 11704 28264 11716
rect 28316 11704 28322 11756
rect 26145 11679 26203 11685
rect 26145 11645 26157 11679
rect 26191 11645 26203 11679
rect 26145 11639 26203 11645
rect 22554 11540 22560 11552
rect 21232 11512 22094 11540
rect 22515 11512 22560 11540
rect 21232 11500 21238 11512
rect 22554 11500 22560 11512
rect 22612 11500 22618 11552
rect 23566 11500 23572 11552
rect 23624 11540 23630 11552
rect 24121 11543 24179 11549
rect 24121 11540 24133 11543
rect 23624 11512 24133 11540
rect 23624 11500 23630 11512
rect 24121 11509 24133 11512
rect 24167 11509 24179 11543
rect 24121 11503 24179 11509
rect 25038 11500 25044 11552
rect 25096 11540 25102 11552
rect 25593 11543 25651 11549
rect 25593 11540 25605 11543
rect 25096 11512 25605 11540
rect 25096 11500 25102 11512
rect 25593 11509 25605 11512
rect 25639 11509 25651 11543
rect 25593 11503 25651 11509
rect 1104 11450 28888 11472
rect 1104 11398 5582 11450
rect 5634 11398 5646 11450
rect 5698 11398 5710 11450
rect 5762 11398 5774 11450
rect 5826 11398 5838 11450
rect 5890 11398 14846 11450
rect 14898 11398 14910 11450
rect 14962 11398 14974 11450
rect 15026 11398 15038 11450
rect 15090 11398 15102 11450
rect 15154 11398 24110 11450
rect 24162 11398 24174 11450
rect 24226 11398 24238 11450
rect 24290 11398 24302 11450
rect 24354 11398 24366 11450
rect 24418 11398 28888 11450
rect 1104 11376 28888 11398
rect 4522 11336 4528 11348
rect 4483 11308 4528 11336
rect 4522 11296 4528 11308
rect 4580 11296 4586 11348
rect 6546 11296 6552 11348
rect 6604 11336 6610 11348
rect 6825 11339 6883 11345
rect 6825 11336 6837 11339
rect 6604 11308 6837 11336
rect 6604 11296 6610 11308
rect 6825 11305 6837 11308
rect 6871 11305 6883 11339
rect 6825 11299 6883 11305
rect 7006 11296 7012 11348
rect 7064 11336 7070 11348
rect 7285 11339 7343 11345
rect 7064 11308 7236 11336
rect 7064 11296 7070 11308
rect 7208 11268 7236 11308
rect 7285 11305 7297 11339
rect 7331 11336 7343 11339
rect 8573 11339 8631 11345
rect 7331 11308 8524 11336
rect 7331 11305 7343 11308
rect 7285 11299 7343 11305
rect 7650 11268 7656 11280
rect 7208 11240 7328 11268
rect 7611 11240 7656 11268
rect 7009 11203 7067 11209
rect 7009 11169 7021 11203
rect 7055 11200 7067 11203
rect 7190 11200 7196 11212
rect 7055 11172 7196 11200
rect 7055 11169 7067 11172
rect 7009 11163 7067 11169
rect 7190 11160 7196 11172
rect 7248 11160 7254 11212
rect 7300 11200 7328 11240
rect 7650 11228 7656 11240
rect 7708 11228 7714 11280
rect 8496 11268 8524 11308
rect 8573 11305 8585 11339
rect 8619 11336 8631 11339
rect 9306 11336 9312 11348
rect 8619 11308 9312 11336
rect 8619 11305 8631 11308
rect 8573 11299 8631 11305
rect 9306 11296 9312 11308
rect 9364 11296 9370 11348
rect 9631 11339 9689 11345
rect 9631 11305 9643 11339
rect 9677 11336 9689 11339
rect 9766 11336 9772 11348
rect 9677 11308 9772 11336
rect 9677 11305 9689 11308
rect 9631 11299 9689 11305
rect 9766 11296 9772 11308
rect 9824 11296 9830 11348
rect 9861 11339 9919 11345
rect 9861 11305 9873 11339
rect 9907 11336 9919 11339
rect 10410 11336 10416 11348
rect 9907 11308 10416 11336
rect 9907 11305 9919 11308
rect 9861 11299 9919 11305
rect 10410 11296 10416 11308
rect 10468 11296 10474 11348
rect 12529 11339 12587 11345
rect 12529 11336 12541 11339
rect 10520 11308 12541 11336
rect 10520 11268 10548 11308
rect 12529 11305 12541 11308
rect 12575 11305 12587 11339
rect 12529 11299 12587 11305
rect 12621 11339 12679 11345
rect 12621 11305 12633 11339
rect 12667 11336 12679 11339
rect 12802 11336 12808 11348
rect 12667 11308 12808 11336
rect 12667 11305 12679 11308
rect 12621 11299 12679 11305
rect 12802 11296 12808 11308
rect 12860 11296 12866 11348
rect 15105 11339 15163 11345
rect 15105 11305 15117 11339
rect 15151 11336 15163 11339
rect 15470 11336 15476 11348
rect 15151 11308 15476 11336
rect 15151 11305 15163 11308
rect 15105 11299 15163 11305
rect 15470 11296 15476 11308
rect 15528 11296 15534 11348
rect 15654 11296 15660 11348
rect 15712 11336 15718 11348
rect 15749 11339 15807 11345
rect 15749 11336 15761 11339
rect 15712 11308 15761 11336
rect 15712 11296 15718 11308
rect 15749 11305 15761 11308
rect 15795 11305 15807 11339
rect 17034 11336 17040 11348
rect 16995 11308 17040 11336
rect 15749 11299 15807 11305
rect 17034 11296 17040 11308
rect 17092 11296 17098 11348
rect 17494 11296 17500 11348
rect 17552 11336 17558 11348
rect 19337 11339 19395 11345
rect 19337 11336 19349 11339
rect 17552 11308 19349 11336
rect 17552 11296 17558 11308
rect 19337 11305 19349 11308
rect 19383 11336 19395 11339
rect 20806 11336 20812 11348
rect 19383 11308 20812 11336
rect 19383 11305 19395 11308
rect 19337 11299 19395 11305
rect 20806 11296 20812 11308
rect 20864 11296 20870 11348
rect 20990 11336 20996 11348
rect 20951 11308 20996 11336
rect 20990 11296 20996 11308
rect 21048 11296 21054 11348
rect 22094 11296 22100 11348
rect 22152 11336 22158 11348
rect 24397 11339 24455 11345
rect 24397 11336 24409 11339
rect 22152 11308 24409 11336
rect 22152 11296 22158 11308
rect 24397 11305 24409 11308
rect 24443 11305 24455 11339
rect 24397 11299 24455 11305
rect 25501 11339 25559 11345
rect 25501 11305 25513 11339
rect 25547 11336 25559 11339
rect 26510 11336 26516 11348
rect 25547 11308 26516 11336
rect 25547 11305 25559 11308
rect 25501 11299 25559 11305
rect 26510 11296 26516 11308
rect 26568 11296 26574 11348
rect 8496 11240 10548 11268
rect 10686 11228 10692 11280
rect 10744 11268 10750 11280
rect 12437 11271 12495 11277
rect 10744 11240 12388 11268
rect 10744 11228 10750 11240
rect 11793 11203 11851 11209
rect 11793 11200 11805 11203
rect 7300 11172 7604 11200
rect 5902 11132 5908 11144
rect 5863 11104 5908 11132
rect 5902 11092 5908 11104
rect 5960 11132 5966 11144
rect 5960 11104 7052 11132
rect 5960 11092 5966 11104
rect 5534 11024 5540 11076
rect 5592 11064 5598 11076
rect 5638 11067 5696 11073
rect 5638 11064 5650 11067
rect 5592 11036 5650 11064
rect 5592 11024 5598 11036
rect 5638 11033 5650 11036
rect 5684 11033 5696 11067
rect 6822 11064 6828 11076
rect 6783 11036 6828 11064
rect 5638 11027 5696 11033
rect 6822 11024 6828 11036
rect 6880 11024 6886 11076
rect 7024 11064 7052 11104
rect 7098 11092 7104 11144
rect 7156 11132 7162 11144
rect 7576 11141 7604 11172
rect 7760 11172 9076 11200
rect 7760 11144 7788 11172
rect 7561 11135 7619 11141
rect 7156 11104 7201 11132
rect 7156 11092 7162 11104
rect 7561 11101 7573 11135
rect 7607 11101 7619 11135
rect 7742 11132 7748 11144
rect 7703 11104 7748 11132
rect 7561 11095 7619 11101
rect 7742 11092 7748 11104
rect 7800 11092 7806 11144
rect 8110 11132 8116 11144
rect 8071 11104 8116 11132
rect 8110 11092 8116 11104
rect 8168 11092 8174 11144
rect 8202 11092 8208 11144
rect 8260 11132 8266 11144
rect 8389 11135 8447 11141
rect 8260 11104 8305 11132
rect 8260 11092 8266 11104
rect 8389 11101 8401 11135
rect 8435 11132 8447 11135
rect 8846 11132 8852 11144
rect 8435 11104 8852 11132
rect 8435 11101 8447 11104
rect 8389 11095 8447 11101
rect 8846 11092 8852 11104
rect 8904 11092 8910 11144
rect 8294 11064 8300 11076
rect 7024 11036 8300 11064
rect 8294 11024 8300 11036
rect 8352 11064 8358 11076
rect 8938 11064 8944 11076
rect 8352 11036 8944 11064
rect 8352 11024 8358 11036
rect 8938 11024 8944 11036
rect 8996 11024 9002 11076
rect 9048 11064 9076 11172
rect 9140 11172 11805 11200
rect 9140 11141 9168 11172
rect 11793 11169 11805 11172
rect 11839 11200 11851 11203
rect 12066 11200 12072 11212
rect 11839 11172 12072 11200
rect 11839 11169 11851 11172
rect 11793 11163 11851 11169
rect 12066 11160 12072 11172
rect 12124 11160 12130 11212
rect 9125 11135 9183 11141
rect 9125 11101 9137 11135
rect 9171 11101 9183 11135
rect 9490 11132 9496 11144
rect 9451 11104 9496 11132
rect 9125 11095 9183 11101
rect 9490 11092 9496 11104
rect 9548 11092 9554 11144
rect 9769 11135 9827 11141
rect 9769 11101 9781 11135
rect 9815 11132 9827 11135
rect 9858 11132 9864 11144
rect 9815 11104 9864 11132
rect 9815 11101 9827 11104
rect 9769 11095 9827 11101
rect 9858 11092 9864 11104
rect 9916 11092 9922 11144
rect 9953 11135 10011 11141
rect 9953 11101 9965 11135
rect 9999 11132 10011 11135
rect 10594 11132 10600 11144
rect 9999 11104 10033 11132
rect 10555 11104 10600 11132
rect 9999 11101 10011 11104
rect 9953 11095 10011 11101
rect 9968 11064 9996 11095
rect 10594 11092 10600 11104
rect 10652 11092 10658 11144
rect 10778 11132 10784 11144
rect 10739 11104 10784 11132
rect 10778 11092 10784 11104
rect 10836 11092 10842 11144
rect 10873 11135 10931 11141
rect 10873 11101 10885 11135
rect 10919 11101 10931 11135
rect 10873 11095 10931 11101
rect 10134 11064 10140 11076
rect 9048 11036 10140 11064
rect 10134 11024 10140 11036
rect 10192 11024 10198 11076
rect 10778 10956 10784 11008
rect 10836 10996 10842 11008
rect 10888 10996 10916 11095
rect 10962 11092 10968 11144
rect 11020 11132 11026 11144
rect 12360 11141 12388 11240
rect 12437 11237 12449 11271
rect 12483 11268 12495 11271
rect 13633 11271 13691 11277
rect 13633 11268 13645 11271
rect 12483 11240 13645 11268
rect 12483 11237 12495 11240
rect 12437 11231 12495 11237
rect 13633 11237 13645 11240
rect 13679 11237 13691 11271
rect 14366 11268 14372 11280
rect 14327 11240 14372 11268
rect 13633 11231 13691 11237
rect 14366 11228 14372 11240
rect 14424 11228 14430 11280
rect 14550 11228 14556 11280
rect 14608 11268 14614 11280
rect 14737 11271 14795 11277
rect 14737 11268 14749 11271
rect 14608 11240 14749 11268
rect 14608 11228 14614 11240
rect 14737 11237 14749 11240
rect 14783 11237 14795 11271
rect 14737 11231 14795 11237
rect 16298 11228 16304 11280
rect 16356 11268 16362 11280
rect 16485 11271 16543 11277
rect 16485 11268 16497 11271
rect 16356 11240 16497 11268
rect 16356 11228 16362 11240
rect 16485 11237 16497 11240
rect 16531 11268 16543 11271
rect 16850 11268 16856 11280
rect 16531 11240 16856 11268
rect 16531 11237 16543 11240
rect 16485 11231 16543 11237
rect 16850 11228 16856 11240
rect 16908 11228 16914 11280
rect 23845 11271 23903 11277
rect 23845 11237 23857 11271
rect 23891 11268 23903 11271
rect 24026 11268 24032 11280
rect 23891 11240 24032 11268
rect 23891 11237 23903 11240
rect 23845 11231 23903 11237
rect 24026 11228 24032 11240
rect 24084 11228 24090 11280
rect 27157 11271 27215 11277
rect 27157 11237 27169 11271
rect 27203 11237 27215 11271
rect 27157 11231 27215 11237
rect 15010 11200 15016 11212
rect 14971 11172 15016 11200
rect 15010 11160 15016 11172
rect 15068 11160 15074 11212
rect 15194 11160 15200 11212
rect 15252 11200 15258 11212
rect 15654 11200 15660 11212
rect 15252 11172 15660 11200
rect 15252 11160 15258 11172
rect 15654 11160 15660 11172
rect 15712 11160 15718 11212
rect 23293 11203 23351 11209
rect 23293 11169 23305 11203
rect 23339 11169 23351 11203
rect 23293 11163 23351 11169
rect 23385 11203 23443 11209
rect 23385 11169 23397 11203
rect 23431 11200 23443 11203
rect 23566 11200 23572 11212
rect 23431 11172 23572 11200
rect 23431 11169 23443 11172
rect 23385 11163 23443 11169
rect 12345 11135 12403 11141
rect 11020 11104 11065 11132
rect 11020 11092 11026 11104
rect 12345 11101 12357 11135
rect 12391 11101 12403 11135
rect 12345 11095 12403 11101
rect 12805 11135 12863 11141
rect 12805 11101 12817 11135
rect 12851 11132 12863 11135
rect 12894 11132 12900 11144
rect 12851 11104 12900 11132
rect 12851 11101 12863 11104
rect 12805 11095 12863 11101
rect 12894 11092 12900 11104
rect 12952 11092 12958 11144
rect 13078 11132 13084 11144
rect 13039 11104 13084 11132
rect 13078 11092 13084 11104
rect 13136 11092 13142 11144
rect 13262 11132 13268 11144
rect 13223 11104 13268 11132
rect 13262 11092 13268 11104
rect 13320 11092 13326 11144
rect 13446 11132 13452 11144
rect 13407 11104 13452 11132
rect 13446 11092 13452 11104
rect 13504 11092 13510 11144
rect 14274 11092 14280 11144
rect 14332 11132 14338 11144
rect 14642 11132 14648 11144
rect 14332 11104 14648 11132
rect 14332 11092 14338 11104
rect 14642 11092 14648 11104
rect 14700 11132 14706 11144
rect 14921 11135 14979 11141
rect 14921 11132 14933 11135
rect 14700 11104 14933 11132
rect 14700 11092 14706 11104
rect 14921 11101 14933 11104
rect 14967 11101 14979 11135
rect 15028 11132 15056 11160
rect 16669 11135 16727 11141
rect 16669 11132 16681 11135
rect 15028 11104 16681 11132
rect 14921 11095 14979 11101
rect 16669 11101 16681 11104
rect 16715 11101 16727 11135
rect 16669 11095 16727 11101
rect 11146 11024 11152 11076
rect 11204 11064 11210 11076
rect 11609 11067 11667 11073
rect 11609 11064 11621 11067
rect 11204 11036 11621 11064
rect 11204 11024 11210 11036
rect 11609 11033 11621 11036
rect 11655 11064 11667 11067
rect 12986 11064 12992 11076
rect 11655 11036 12992 11064
rect 11655 11033 11667 11036
rect 11609 11027 11667 11033
rect 12986 11024 12992 11036
rect 13044 11024 13050 11076
rect 13354 11024 13360 11076
rect 13412 11064 13418 11076
rect 13412 11036 13457 11064
rect 13412 11024 13418 11036
rect 13906 11024 13912 11076
rect 13964 11064 13970 11076
rect 14185 11067 14243 11073
rect 14185 11064 14197 11067
rect 13964 11036 14197 11064
rect 13964 11024 13970 11036
rect 14185 11033 14197 11036
rect 14231 11033 14243 11067
rect 15194 11064 15200 11076
rect 15155 11036 15200 11064
rect 14185 11027 14243 11033
rect 15194 11024 15200 11036
rect 15252 11024 15258 11076
rect 16114 11064 16120 11076
rect 16075 11036 16120 11064
rect 16114 11024 16120 11036
rect 16172 11024 16178 11076
rect 11238 10996 11244 11008
rect 10836 10968 10916 10996
rect 11199 10968 11244 10996
rect 10836 10956 10842 10968
rect 11238 10956 11244 10968
rect 11296 10956 11302 11008
rect 12066 10996 12072 11008
rect 12027 10968 12072 10996
rect 12066 10956 12072 10968
rect 12124 10956 12130 11008
rect 16684 10996 16712 11095
rect 18046 11092 18052 11144
rect 18104 11132 18110 11144
rect 18785 11135 18843 11141
rect 18785 11132 18797 11135
rect 18104 11104 18797 11132
rect 18104 11092 18110 11104
rect 18785 11101 18797 11104
rect 18831 11132 18843 11135
rect 19242 11132 19248 11144
rect 18831 11104 19248 11132
rect 18831 11101 18843 11104
rect 18785 11095 18843 11101
rect 19242 11092 19248 11104
rect 19300 11132 19306 11144
rect 19613 11135 19671 11141
rect 19613 11132 19625 11135
rect 19300 11104 19625 11132
rect 19300 11092 19306 11104
rect 19613 11101 19625 11104
rect 19659 11132 19671 11135
rect 21361 11135 21419 11141
rect 21361 11132 21373 11135
rect 19659 11104 21373 11132
rect 19659 11101 19671 11104
rect 19613 11095 19671 11101
rect 20088 11076 20116 11104
rect 21361 11101 21373 11104
rect 21407 11101 21419 11135
rect 23308 11132 23336 11163
rect 23566 11160 23572 11172
rect 23624 11160 23630 11212
rect 24857 11203 24915 11209
rect 24857 11169 24869 11203
rect 24903 11169 24915 11203
rect 25038 11200 25044 11212
rect 24999 11172 25044 11200
rect 24857 11163 24915 11169
rect 24872 11132 24900 11163
rect 25038 11160 25044 11172
rect 25096 11160 25102 11212
rect 24946 11132 24952 11144
rect 23308 11104 24952 11132
rect 21361 11095 21419 11101
rect 24946 11092 24952 11104
rect 25004 11092 25010 11144
rect 25130 11132 25136 11144
rect 25091 11104 25136 11132
rect 25130 11092 25136 11104
rect 25188 11092 25194 11144
rect 25774 11132 25780 11144
rect 25735 11104 25780 11132
rect 25774 11092 25780 11104
rect 25832 11092 25838 11144
rect 26326 11092 26332 11144
rect 26384 11132 26390 11144
rect 27172 11132 27200 11231
rect 26384 11104 27200 11132
rect 26384 11092 26390 11104
rect 17770 11024 17776 11076
rect 17828 11064 17834 11076
rect 18518 11067 18576 11073
rect 18518 11064 18530 11067
rect 17828 11036 18530 11064
rect 17828 11024 17834 11036
rect 18518 11033 18530 11036
rect 18564 11033 18576 11067
rect 18518 11027 18576 11033
rect 18966 11024 18972 11076
rect 19024 11064 19030 11076
rect 19858 11067 19916 11073
rect 19858 11064 19870 11067
rect 19024 11036 19870 11064
rect 19024 11024 19030 11036
rect 19858 11033 19870 11036
rect 19904 11033 19916 11067
rect 19858 11027 19916 11033
rect 20070 11024 20076 11076
rect 20128 11024 20134 11076
rect 21628 11067 21686 11073
rect 21628 11033 21640 11067
rect 21674 11064 21686 11067
rect 22554 11064 22560 11076
rect 21674 11036 22560 11064
rect 21674 11033 21686 11036
rect 21628 11027 21686 11033
rect 22554 11024 22560 11036
rect 22612 11024 22618 11076
rect 23477 11067 23535 11073
rect 23477 11064 23489 11067
rect 22756 11036 23489 11064
rect 17405 10999 17463 11005
rect 17405 10996 17417 10999
rect 16684 10968 17417 10996
rect 17405 10965 17417 10968
rect 17451 10965 17463 10999
rect 17405 10959 17463 10965
rect 22462 10956 22468 11008
rect 22520 10996 22526 11008
rect 22756 11005 22784 11036
rect 23477 11033 23489 11036
rect 23523 11033 23535 11067
rect 23477 11027 23535 11033
rect 26044 11067 26102 11073
rect 26044 11033 26056 11067
rect 26090 11064 26102 11067
rect 26418 11064 26424 11076
rect 26090 11036 26424 11064
rect 26090 11033 26102 11036
rect 26044 11027 26102 11033
rect 26418 11024 26424 11036
rect 26476 11024 26482 11076
rect 22741 10999 22799 11005
rect 22741 10996 22753 10999
rect 22520 10968 22753 10996
rect 22520 10956 22526 10968
rect 22741 10965 22753 10968
rect 22787 10965 22799 10999
rect 22741 10959 22799 10965
rect 1104 10906 28888 10928
rect 1104 10854 10214 10906
rect 10266 10854 10278 10906
rect 10330 10854 10342 10906
rect 10394 10854 10406 10906
rect 10458 10854 10470 10906
rect 10522 10854 19478 10906
rect 19530 10854 19542 10906
rect 19594 10854 19606 10906
rect 19658 10854 19670 10906
rect 19722 10854 19734 10906
rect 19786 10854 28888 10906
rect 1104 10832 28888 10854
rect 7834 10792 7840 10804
rect 7795 10764 7840 10792
rect 7834 10752 7840 10764
rect 7892 10792 7898 10804
rect 8110 10792 8116 10804
rect 7892 10764 8116 10792
rect 7892 10752 7898 10764
rect 8110 10752 8116 10764
rect 8168 10752 8174 10804
rect 8849 10795 8907 10801
rect 8849 10761 8861 10795
rect 8895 10761 8907 10795
rect 10870 10792 10876 10804
rect 10831 10764 10876 10792
rect 8849 10755 8907 10761
rect 7190 10724 7196 10736
rect 6840 10696 7196 10724
rect 5629 10659 5687 10665
rect 5629 10625 5641 10659
rect 5675 10656 5687 10659
rect 5994 10656 6000 10668
rect 5675 10628 6000 10656
rect 5675 10625 5687 10628
rect 5629 10619 5687 10625
rect 5994 10616 6000 10628
rect 6052 10616 6058 10668
rect 6840 10665 6868 10696
rect 7190 10684 7196 10696
rect 7248 10684 7254 10736
rect 8864 10724 8892 10755
rect 10870 10752 10876 10764
rect 10928 10752 10934 10804
rect 10962 10752 10968 10804
rect 11020 10792 11026 10804
rect 11020 10764 12434 10792
rect 11020 10752 11026 10764
rect 9370 10727 9428 10733
rect 9370 10724 9382 10727
rect 8864 10696 9382 10724
rect 9370 10693 9382 10696
rect 9416 10693 9428 10727
rect 9370 10687 9428 10693
rect 9674 10684 9680 10736
rect 9732 10724 9738 10736
rect 10980 10724 11008 10752
rect 9732 10696 11008 10724
rect 9732 10684 9738 10696
rect 6641 10659 6699 10665
rect 6641 10625 6653 10659
rect 6687 10625 6699 10659
rect 6641 10619 6699 10625
rect 6825 10659 6883 10665
rect 6825 10625 6837 10659
rect 6871 10625 6883 10659
rect 7098 10656 7104 10668
rect 7059 10628 7104 10656
rect 6825 10619 6883 10625
rect 6656 10588 6684 10619
rect 7098 10616 7104 10628
rect 7156 10616 7162 10668
rect 7377 10659 7435 10665
rect 7377 10625 7389 10659
rect 7423 10656 7435 10659
rect 7466 10656 7472 10668
rect 7423 10628 7472 10656
rect 7423 10625 7435 10628
rect 7377 10619 7435 10625
rect 7466 10616 7472 10628
rect 7524 10616 7530 10668
rect 7742 10656 7748 10668
rect 7703 10628 7748 10656
rect 7742 10616 7748 10628
rect 7800 10616 7806 10668
rect 8662 10656 8668 10668
rect 8623 10628 8668 10656
rect 8662 10616 8668 10628
rect 8720 10616 8726 10668
rect 8938 10616 8944 10668
rect 8996 10656 9002 10668
rect 9125 10659 9183 10665
rect 9125 10656 9137 10659
rect 8996 10628 9137 10656
rect 8996 10616 9002 10628
rect 9125 10625 9137 10628
rect 9171 10625 9183 10659
rect 9125 10619 9183 10625
rect 10134 10616 10140 10668
rect 10192 10656 10198 10668
rect 10980 10665 11008 10696
rect 11238 10684 11244 10736
rect 11296 10724 11302 10736
rect 11762 10727 11820 10733
rect 11762 10724 11774 10727
rect 11296 10696 11774 10724
rect 11296 10684 11302 10696
rect 11762 10693 11774 10696
rect 11808 10693 11820 10727
rect 11762 10687 11820 10693
rect 11974 10684 11980 10736
rect 12032 10684 12038 10736
rect 10781 10659 10839 10665
rect 10781 10656 10793 10659
rect 10192 10628 10793 10656
rect 10192 10616 10198 10628
rect 10781 10625 10793 10628
rect 10827 10625 10839 10659
rect 10781 10619 10839 10625
rect 10965 10659 11023 10665
rect 10965 10625 10977 10659
rect 11011 10625 11023 10659
rect 10965 10619 11023 10625
rect 11517 10659 11575 10665
rect 11517 10625 11529 10659
rect 11563 10656 11575 10659
rect 11992 10656 12020 10684
rect 11563 10628 12020 10656
rect 12406 10656 12434 10764
rect 14182 10752 14188 10804
rect 14240 10792 14246 10804
rect 16666 10792 16672 10804
rect 14240 10764 16672 10792
rect 14240 10752 14246 10764
rect 16666 10752 16672 10764
rect 16724 10792 16730 10804
rect 16945 10795 17003 10801
rect 16945 10792 16957 10795
rect 16724 10764 16957 10792
rect 16724 10752 16730 10764
rect 16945 10761 16957 10764
rect 16991 10761 17003 10795
rect 17497 10795 17555 10801
rect 17497 10792 17509 10795
rect 16945 10755 17003 10761
rect 17052 10764 17509 10792
rect 14366 10684 14372 10736
rect 14424 10724 14430 10736
rect 17052 10733 17080 10764
rect 17497 10761 17509 10764
rect 17543 10761 17555 10795
rect 19242 10792 19248 10804
rect 19203 10764 19248 10792
rect 17497 10755 17555 10761
rect 19242 10752 19248 10764
rect 19300 10752 19306 10804
rect 20254 10752 20260 10804
rect 20312 10792 20318 10804
rect 20717 10795 20775 10801
rect 20717 10792 20729 10795
rect 20312 10764 20729 10792
rect 20312 10752 20318 10764
rect 20717 10761 20729 10764
rect 20763 10761 20775 10795
rect 20717 10755 20775 10761
rect 20990 10752 20996 10804
rect 21048 10792 21054 10804
rect 25777 10795 25835 10801
rect 25777 10792 25789 10795
rect 21048 10764 25789 10792
rect 21048 10752 21054 10764
rect 25777 10761 25789 10764
rect 25823 10761 25835 10795
rect 26418 10792 26424 10804
rect 26379 10764 26424 10792
rect 25777 10755 25835 10761
rect 26418 10752 26424 10764
rect 26476 10752 26482 10804
rect 14461 10727 14519 10733
rect 14461 10724 14473 10727
rect 14424 10696 14473 10724
rect 14424 10684 14430 10696
rect 14461 10693 14473 10696
rect 14507 10693 14519 10727
rect 14461 10687 14519 10693
rect 14645 10727 14703 10733
rect 14645 10693 14657 10727
rect 14691 10724 14703 10727
rect 15013 10727 15071 10733
rect 15013 10724 15025 10727
rect 14691 10696 15025 10724
rect 14691 10693 14703 10696
rect 14645 10687 14703 10693
rect 15013 10693 15025 10696
rect 15059 10724 15071 10727
rect 17037 10727 17095 10733
rect 17037 10724 17049 10727
rect 15059 10696 17049 10724
rect 15059 10693 15071 10696
rect 15013 10687 15071 10693
rect 17037 10693 17049 10696
rect 17083 10693 17095 10727
rect 17037 10687 17095 10693
rect 18322 10684 18328 10736
rect 18380 10724 18386 10736
rect 18610 10727 18668 10733
rect 18610 10724 18622 10727
rect 18380 10696 18622 10724
rect 18380 10684 18386 10696
rect 18610 10693 18622 10696
rect 18656 10693 18668 10727
rect 18610 10687 18668 10693
rect 13262 10656 13268 10668
rect 12406 10628 13268 10656
rect 11563 10625 11575 10628
rect 11517 10619 11575 10625
rect 13262 10616 13268 10628
rect 13320 10656 13326 10668
rect 13449 10659 13507 10665
rect 13449 10656 13461 10659
rect 13320 10628 13461 10656
rect 13320 10616 13326 10628
rect 13449 10625 13461 10628
rect 13495 10625 13507 10659
rect 15286 10656 15292 10668
rect 15247 10628 15292 10656
rect 13449 10619 13507 10625
rect 15286 10616 15292 10628
rect 15344 10616 15350 10668
rect 18877 10659 18935 10665
rect 18877 10625 18889 10659
rect 18923 10656 18935 10659
rect 19260 10656 19288 10752
rect 19337 10727 19395 10733
rect 19337 10693 19349 10727
rect 19383 10724 19395 10727
rect 21174 10724 21180 10736
rect 19383 10696 21180 10724
rect 19383 10693 19395 10696
rect 19337 10687 19395 10693
rect 21174 10684 21180 10696
rect 21232 10684 21238 10736
rect 21358 10724 21364 10736
rect 21319 10696 21364 10724
rect 21358 10684 21364 10696
rect 21416 10684 21422 10736
rect 22462 10724 22468 10736
rect 22423 10696 22468 10724
rect 22462 10684 22468 10696
rect 22520 10684 22526 10736
rect 23744 10727 23802 10733
rect 23744 10693 23756 10727
rect 23790 10724 23802 10727
rect 23842 10724 23848 10736
rect 23790 10696 23848 10724
rect 23790 10693 23802 10696
rect 23744 10687 23802 10693
rect 23842 10684 23848 10696
rect 23900 10684 23906 10736
rect 19886 10656 19892 10668
rect 18923 10628 19288 10656
rect 19799 10628 19892 10656
rect 18923 10625 18935 10628
rect 18877 10619 18935 10625
rect 19886 10616 19892 10628
rect 19944 10616 19950 10668
rect 20070 10656 20076 10668
rect 20031 10628 20076 10656
rect 20070 10616 20076 10628
rect 20128 10616 20134 10668
rect 20346 10656 20352 10668
rect 20307 10628 20352 10656
rect 20346 10616 20352 10628
rect 20404 10616 20410 10668
rect 20533 10659 20591 10665
rect 20533 10625 20545 10659
rect 20579 10625 20591 10659
rect 20533 10619 20591 10625
rect 7760 10588 7788 10616
rect 13173 10591 13231 10597
rect 13173 10588 13185 10591
rect 6656 10560 7788 10588
rect 12912 10560 13185 10588
rect 6914 10480 6920 10532
rect 6972 10520 6978 10532
rect 7377 10523 7435 10529
rect 7377 10520 7389 10523
rect 6972 10492 7389 10520
rect 6972 10480 6978 10492
rect 7377 10489 7389 10492
rect 7423 10489 7435 10523
rect 7377 10483 7435 10489
rect 12802 10480 12808 10532
rect 12860 10520 12866 10532
rect 12912 10529 12940 10560
rect 13173 10557 13185 10560
rect 13219 10557 13231 10591
rect 13173 10551 13231 10557
rect 13906 10548 13912 10600
rect 13964 10588 13970 10600
rect 15197 10591 15255 10597
rect 15197 10588 15209 10591
rect 13964 10560 15209 10588
rect 13964 10548 13970 10560
rect 15197 10557 15209 10560
rect 15243 10557 15255 10591
rect 19904 10588 19932 10616
rect 20548 10588 20576 10619
rect 20898 10616 20904 10668
rect 20956 10656 20962 10668
rect 20993 10659 21051 10665
rect 20993 10656 21005 10659
rect 20956 10628 21005 10656
rect 20956 10616 20962 10628
rect 20993 10625 21005 10628
rect 21039 10625 21051 10659
rect 20993 10619 21051 10625
rect 21450 10616 21456 10668
rect 21508 10656 21514 10668
rect 22373 10659 22431 10665
rect 22373 10656 22385 10659
rect 21508 10628 22385 10656
rect 21508 10616 21514 10628
rect 22373 10625 22385 10628
rect 22419 10625 22431 10659
rect 22373 10619 22431 10625
rect 23201 10659 23259 10665
rect 23201 10625 23213 10659
rect 23247 10625 23259 10659
rect 23474 10656 23480 10668
rect 23435 10628 23480 10656
rect 23201 10619 23259 10625
rect 22554 10588 22560 10600
rect 15197 10551 15255 10557
rect 19260 10560 20576 10588
rect 22515 10560 22560 10588
rect 12897 10523 12955 10529
rect 12897 10520 12909 10523
rect 12860 10492 12909 10520
rect 12860 10480 12866 10492
rect 12897 10489 12909 10492
rect 12943 10489 12955 10523
rect 12897 10483 12955 10489
rect 13538 10480 13544 10532
rect 13596 10520 13602 10532
rect 13596 10492 18000 10520
rect 13596 10480 13602 10492
rect 1394 10452 1400 10464
rect 1355 10424 1400 10452
rect 1394 10412 1400 10424
rect 1452 10412 1458 10464
rect 5442 10452 5448 10464
rect 5403 10424 5448 10452
rect 5442 10412 5448 10424
rect 5500 10412 5506 10464
rect 6822 10452 6828 10464
rect 6783 10424 6828 10452
rect 6822 10412 6828 10424
rect 6880 10412 6886 10464
rect 7098 10412 7104 10464
rect 7156 10452 7162 10464
rect 7558 10452 7564 10464
rect 7156 10424 7564 10452
rect 7156 10412 7162 10424
rect 7558 10412 7564 10424
rect 7616 10452 7622 10464
rect 8297 10455 8355 10461
rect 8297 10452 8309 10455
rect 7616 10424 8309 10452
rect 7616 10412 7622 10424
rect 8297 10421 8309 10424
rect 8343 10452 8355 10455
rect 9030 10452 9036 10464
rect 8343 10424 9036 10452
rect 8343 10421 8355 10424
rect 8297 10415 8355 10421
rect 9030 10412 9036 10424
rect 9088 10412 9094 10464
rect 10505 10455 10563 10461
rect 10505 10421 10517 10455
rect 10551 10452 10563 10455
rect 11146 10452 11152 10464
rect 10551 10424 11152 10452
rect 10551 10421 10563 10424
rect 10505 10415 10563 10421
rect 11146 10412 11152 10424
rect 11204 10412 11210 10464
rect 14090 10412 14096 10464
rect 14148 10452 14154 10464
rect 14277 10455 14335 10461
rect 14277 10452 14289 10455
rect 14148 10424 14289 10452
rect 14148 10412 14154 10424
rect 14277 10421 14289 10424
rect 14323 10421 14335 10455
rect 14277 10415 14335 10421
rect 14458 10412 14464 10464
rect 14516 10452 14522 10464
rect 15013 10455 15071 10461
rect 15013 10452 15025 10455
rect 14516 10424 15025 10452
rect 14516 10412 14522 10424
rect 15013 10421 15025 10424
rect 15059 10421 15071 10455
rect 15013 10415 15071 10421
rect 15194 10412 15200 10464
rect 15252 10452 15258 10464
rect 15473 10455 15531 10461
rect 15473 10452 15485 10455
rect 15252 10424 15485 10452
rect 15252 10412 15258 10424
rect 15473 10421 15485 10424
rect 15519 10452 15531 10455
rect 15838 10452 15844 10464
rect 15519 10424 15844 10452
rect 15519 10421 15531 10424
rect 15473 10415 15531 10421
rect 15838 10412 15844 10424
rect 15896 10412 15902 10464
rect 17972 10452 18000 10492
rect 19260 10452 19288 10560
rect 22554 10548 22560 10560
rect 22612 10548 22618 10600
rect 19426 10480 19432 10532
rect 19484 10520 19490 10532
rect 20346 10520 20352 10532
rect 19484 10492 20352 10520
rect 19484 10480 19490 10492
rect 20346 10480 20352 10492
rect 20404 10480 20410 10532
rect 17972 10424 19288 10452
rect 19334 10412 19340 10464
rect 19392 10452 19398 10464
rect 19705 10455 19763 10461
rect 19705 10452 19717 10455
rect 19392 10424 19717 10452
rect 19392 10412 19398 10424
rect 19705 10421 19717 10424
rect 19751 10421 19763 10455
rect 19705 10415 19763 10421
rect 21910 10412 21916 10464
rect 21968 10452 21974 10464
rect 22005 10455 22063 10461
rect 22005 10452 22017 10455
rect 21968 10424 22017 10452
rect 21968 10412 21974 10424
rect 22005 10421 22017 10424
rect 22051 10421 22063 10455
rect 23014 10452 23020 10464
rect 22975 10424 23020 10452
rect 22005 10415 22063 10421
rect 23014 10412 23020 10424
rect 23072 10412 23078 10464
rect 23216 10452 23244 10619
rect 23474 10616 23480 10628
rect 23532 10616 23538 10668
rect 26510 10616 26516 10668
rect 26568 10656 26574 10668
rect 26605 10659 26663 10665
rect 26605 10656 26617 10659
rect 26568 10628 26617 10656
rect 26568 10616 26574 10628
rect 26605 10625 26617 10628
rect 26651 10625 26663 10659
rect 28074 10656 28080 10668
rect 28035 10628 28080 10656
rect 26605 10619 26663 10625
rect 28074 10616 28080 10628
rect 28132 10616 28138 10668
rect 25498 10588 25504 10600
rect 25459 10560 25504 10588
rect 25498 10548 25504 10560
rect 25556 10548 25562 10600
rect 25682 10588 25688 10600
rect 25643 10560 25688 10588
rect 25682 10548 25688 10560
rect 25740 10548 25746 10600
rect 24857 10523 24915 10529
rect 24857 10489 24869 10523
rect 24903 10520 24915 10523
rect 25130 10520 25136 10532
rect 24903 10492 25136 10520
rect 24903 10489 24915 10492
rect 24857 10483 24915 10489
rect 25130 10480 25136 10492
rect 25188 10480 25194 10532
rect 24670 10452 24676 10464
rect 23216 10424 24676 10452
rect 24670 10412 24676 10424
rect 24728 10412 24734 10464
rect 26142 10452 26148 10464
rect 26103 10424 26148 10452
rect 26142 10412 26148 10424
rect 26200 10412 26206 10464
rect 28258 10452 28264 10464
rect 28219 10424 28264 10452
rect 28258 10412 28264 10424
rect 28316 10412 28322 10464
rect 1104 10362 28888 10384
rect 1104 10310 5582 10362
rect 5634 10310 5646 10362
rect 5698 10310 5710 10362
rect 5762 10310 5774 10362
rect 5826 10310 5838 10362
rect 5890 10310 14846 10362
rect 14898 10310 14910 10362
rect 14962 10310 14974 10362
rect 15026 10310 15038 10362
rect 15090 10310 15102 10362
rect 15154 10310 24110 10362
rect 24162 10310 24174 10362
rect 24226 10310 24238 10362
rect 24290 10310 24302 10362
rect 24354 10310 24366 10362
rect 24418 10310 28888 10362
rect 1104 10288 28888 10310
rect 7282 10248 7288 10260
rect 7243 10220 7288 10248
rect 7282 10208 7288 10220
rect 7340 10208 7346 10260
rect 8386 10208 8392 10260
rect 8444 10248 8450 10260
rect 8941 10251 8999 10257
rect 8941 10248 8953 10251
rect 8444 10220 8953 10248
rect 8444 10208 8450 10220
rect 8941 10217 8953 10220
rect 8987 10217 8999 10251
rect 8941 10211 8999 10217
rect 9030 10208 9036 10260
rect 9088 10248 9094 10260
rect 13173 10251 13231 10257
rect 9088 10220 12434 10248
rect 9088 10208 9094 10220
rect 6549 10183 6607 10189
rect 6549 10149 6561 10183
rect 6595 10149 6607 10183
rect 6549 10143 6607 10149
rect 6564 10112 6592 10143
rect 6822 10140 6828 10192
rect 6880 10180 6886 10192
rect 10778 10180 10784 10192
rect 6880 10152 10784 10180
rect 6880 10140 6886 10152
rect 7561 10115 7619 10121
rect 7561 10112 7573 10115
rect 6564 10084 7573 10112
rect 7561 10081 7573 10084
rect 7607 10112 7619 10115
rect 7742 10112 7748 10124
rect 7607 10084 7748 10112
rect 7607 10081 7619 10084
rect 7561 10075 7619 10081
rect 7742 10072 7748 10084
rect 7800 10072 7806 10124
rect 9122 10112 9128 10124
rect 9083 10084 9128 10112
rect 9122 10072 9128 10084
rect 9180 10072 9186 10124
rect 9416 10121 9444 10152
rect 10778 10140 10784 10152
rect 10836 10140 10842 10192
rect 12406 10180 12434 10220
rect 13173 10217 13185 10251
rect 13219 10248 13231 10251
rect 13354 10248 13360 10260
rect 13219 10220 13360 10248
rect 13219 10217 13231 10220
rect 13173 10211 13231 10217
rect 13354 10208 13360 10220
rect 13412 10208 13418 10260
rect 13446 10208 13452 10260
rect 13504 10248 13510 10260
rect 13541 10251 13599 10257
rect 13541 10248 13553 10251
rect 13504 10220 13553 10248
rect 13504 10208 13510 10220
rect 13541 10217 13553 10220
rect 13587 10217 13599 10251
rect 22370 10248 22376 10260
rect 13541 10211 13599 10217
rect 15396 10220 16436 10248
rect 22331 10220 22376 10248
rect 15396 10180 15424 10220
rect 12406 10152 15424 10180
rect 15473 10183 15531 10189
rect 15473 10149 15485 10183
rect 15519 10180 15531 10183
rect 16298 10180 16304 10192
rect 15519 10152 16304 10180
rect 15519 10149 15531 10152
rect 15473 10143 15531 10149
rect 16298 10140 16304 10152
rect 16356 10140 16362 10192
rect 9401 10115 9459 10121
rect 9401 10081 9413 10115
rect 9447 10081 9459 10115
rect 11146 10112 11152 10124
rect 11107 10084 11152 10112
rect 9401 10075 9459 10081
rect 11146 10072 11152 10084
rect 11204 10072 11210 10124
rect 11425 10115 11483 10121
rect 11425 10081 11437 10115
rect 11471 10112 11483 10115
rect 12250 10112 12256 10124
rect 11471 10084 12256 10112
rect 11471 10081 11483 10084
rect 11425 10075 11483 10081
rect 12250 10072 12256 10084
rect 12308 10072 12314 10124
rect 14921 10115 14979 10121
rect 13648 10084 14320 10112
rect 5169 10047 5227 10053
rect 5169 10013 5181 10047
rect 5215 10044 5227 10047
rect 5902 10044 5908 10056
rect 5215 10016 5908 10044
rect 5215 10013 5227 10016
rect 5169 10007 5227 10013
rect 5902 10004 5908 10016
rect 5960 10004 5966 10056
rect 6917 10047 6975 10053
rect 6917 10013 6929 10047
rect 6963 10013 6975 10047
rect 7098 10044 7104 10056
rect 7059 10016 7104 10044
rect 6917 10007 6975 10013
rect 5442 9985 5448 9988
rect 5436 9976 5448 9985
rect 5403 9948 5448 9976
rect 5436 9939 5448 9948
rect 5442 9936 5448 9939
rect 5500 9936 5506 9988
rect 6932 9976 6960 10007
rect 7098 10004 7104 10016
rect 7156 10004 7162 10056
rect 7837 10047 7895 10053
rect 7837 10013 7849 10047
rect 7883 10044 7895 10047
rect 8294 10044 8300 10056
rect 7883 10016 8300 10044
rect 7883 10013 7895 10016
rect 7837 10007 7895 10013
rect 8294 10004 8300 10016
rect 8352 10004 8358 10056
rect 9214 10044 9220 10056
rect 9175 10016 9220 10044
rect 9214 10004 9220 10016
rect 9272 10004 9278 10056
rect 9306 10004 9312 10056
rect 9364 10044 9370 10056
rect 12802 10044 12808 10056
rect 9364 10016 9409 10044
rect 12763 10016 12808 10044
rect 9364 10004 9370 10016
rect 12802 10004 12808 10016
rect 12860 10004 12866 10056
rect 13262 10004 13268 10056
rect 13320 10044 13326 10056
rect 13648 10053 13676 10084
rect 13449 10047 13507 10053
rect 13449 10044 13461 10047
rect 13320 10016 13461 10044
rect 13320 10004 13326 10016
rect 13449 10013 13461 10016
rect 13495 10013 13507 10047
rect 13449 10007 13507 10013
rect 13633 10047 13691 10053
rect 13633 10013 13645 10047
rect 13679 10013 13691 10047
rect 13633 10007 13691 10013
rect 14093 10047 14151 10053
rect 14093 10013 14105 10047
rect 14139 10044 14151 10047
rect 14182 10044 14188 10056
rect 14139 10016 14188 10044
rect 14139 10013 14151 10016
rect 14093 10007 14151 10013
rect 14182 10004 14188 10016
rect 14240 10004 14246 10056
rect 14292 10053 14320 10084
rect 14921 10081 14933 10115
rect 14967 10112 14979 10115
rect 15565 10115 15623 10121
rect 15565 10112 15577 10115
rect 14967 10084 15577 10112
rect 14967 10081 14979 10084
rect 14921 10075 14979 10081
rect 15565 10081 15577 10084
rect 15611 10112 15623 10115
rect 15838 10112 15844 10124
rect 15611 10084 15844 10112
rect 15611 10081 15623 10084
rect 15565 10075 15623 10081
rect 15838 10072 15844 10084
rect 15896 10072 15902 10124
rect 16408 10112 16436 10220
rect 22370 10208 22376 10220
rect 22428 10208 22434 10260
rect 22554 10208 22560 10260
rect 22612 10248 22618 10260
rect 25593 10251 25651 10257
rect 22612 10220 24256 10248
rect 22612 10208 22618 10220
rect 17678 10180 17684 10192
rect 17639 10152 17684 10180
rect 17678 10140 17684 10152
rect 17736 10140 17742 10192
rect 16408 10084 18368 10112
rect 18340 10056 18368 10084
rect 19242 10072 19248 10124
rect 19300 10112 19306 10124
rect 19797 10115 19855 10121
rect 19797 10112 19809 10115
rect 19300 10084 19809 10112
rect 19300 10072 19306 10084
rect 19797 10081 19809 10084
rect 19843 10081 19855 10115
rect 19797 10075 19855 10081
rect 21821 10115 21879 10121
rect 21821 10081 21833 10115
rect 21867 10081 21879 10115
rect 21821 10075 21879 10081
rect 14277 10047 14335 10053
rect 14277 10013 14289 10047
rect 14323 10044 14335 10047
rect 14366 10044 14372 10056
rect 14323 10016 14372 10044
rect 14323 10013 14335 10016
rect 14277 10007 14335 10013
rect 14366 10004 14372 10016
rect 14424 10004 14430 10056
rect 14734 10044 14740 10056
rect 14695 10016 14740 10044
rect 14734 10004 14740 10016
rect 14792 10004 14798 10056
rect 15381 10047 15439 10053
rect 15381 10013 15393 10047
rect 15427 10044 15439 10047
rect 15470 10044 15476 10056
rect 15427 10016 15476 10044
rect 15427 10013 15439 10016
rect 15381 10007 15439 10013
rect 15470 10004 15476 10016
rect 15528 10004 15534 10056
rect 15657 10047 15715 10053
rect 15657 10013 15669 10047
rect 15703 10044 15715 10047
rect 16669 10047 16727 10053
rect 16669 10044 16681 10047
rect 15703 10016 15792 10044
rect 15703 10013 15715 10016
rect 15657 10007 15715 10013
rect 9232 9976 9260 10004
rect 6932 9948 9260 9976
rect 12066 9936 12072 9988
rect 12124 9976 12130 9988
rect 12437 9979 12495 9985
rect 12437 9976 12449 9979
rect 12124 9948 12449 9976
rect 12124 9936 12130 9948
rect 12437 9945 12449 9948
rect 12483 9945 12495 9979
rect 12437 9939 12495 9945
rect 12989 9979 13047 9985
rect 12989 9945 13001 9979
rect 13035 9976 13047 9979
rect 13906 9976 13912 9988
rect 13035 9948 13912 9976
rect 13035 9945 13047 9948
rect 12989 9939 13047 9945
rect 13906 9936 13912 9948
rect 13964 9936 13970 9988
rect 13998 9936 14004 9988
rect 14056 9976 14062 9988
rect 14553 9979 14611 9985
rect 14553 9976 14565 9979
rect 14056 9948 14565 9976
rect 14056 9936 14062 9948
rect 14553 9945 14565 9948
rect 14599 9945 14611 9979
rect 14553 9939 14611 9945
rect 14642 9936 14648 9988
rect 14700 9976 14706 9988
rect 15764 9976 15792 10016
rect 14700 9948 15792 9976
rect 15856 10016 16681 10044
rect 14700 9936 14706 9948
rect 12342 9908 12348 9920
rect 12303 9880 12348 9908
rect 12342 9868 12348 9880
rect 12400 9868 12406 9920
rect 14274 9908 14280 9920
rect 14235 9880 14280 9908
rect 14274 9868 14280 9880
rect 14332 9868 14338 9920
rect 15197 9911 15255 9917
rect 15197 9877 15209 9911
rect 15243 9908 15255 9911
rect 15378 9908 15384 9920
rect 15243 9880 15384 9908
rect 15243 9877 15255 9880
rect 15197 9871 15255 9877
rect 15378 9868 15384 9880
rect 15436 9868 15442 9920
rect 15470 9868 15476 9920
rect 15528 9908 15534 9920
rect 15856 9908 15884 10016
rect 16669 10013 16681 10016
rect 16715 10013 16727 10047
rect 16669 10007 16727 10013
rect 16758 10004 16764 10056
rect 16816 10044 16822 10056
rect 17037 10047 17095 10053
rect 17037 10044 17049 10047
rect 16816 10016 17049 10044
rect 16816 10004 16822 10016
rect 17037 10013 17049 10016
rect 17083 10044 17095 10047
rect 17405 10047 17463 10053
rect 17405 10044 17417 10047
rect 17083 10016 17417 10044
rect 17083 10013 17095 10016
rect 17037 10007 17095 10013
rect 17405 10013 17417 10016
rect 17451 10013 17463 10047
rect 18322 10044 18328 10056
rect 18235 10016 18328 10044
rect 17405 10007 17463 10013
rect 18322 10004 18328 10016
rect 18380 10044 18386 10056
rect 18693 10047 18751 10053
rect 18693 10044 18705 10047
rect 18380 10016 18705 10044
rect 18380 10004 18386 10016
rect 18693 10013 18705 10016
rect 18739 10044 18751 10047
rect 19150 10044 19156 10056
rect 18739 10016 19156 10044
rect 18739 10013 18751 10016
rect 18693 10007 18751 10013
rect 19150 10004 19156 10016
rect 19208 10004 19214 10056
rect 19334 10044 19340 10056
rect 19295 10016 19340 10044
rect 19334 10004 19340 10016
rect 19392 10004 19398 10056
rect 21836 10044 21864 10075
rect 21910 10072 21916 10124
rect 21968 10112 21974 10124
rect 24228 10112 24256 10220
rect 25593 10217 25605 10251
rect 25639 10248 25651 10251
rect 25682 10248 25688 10260
rect 25639 10220 25688 10248
rect 25639 10217 25651 10220
rect 25593 10211 25651 10217
rect 25682 10208 25688 10220
rect 25740 10208 25746 10260
rect 24489 10115 24547 10121
rect 24489 10112 24501 10115
rect 21968 10084 22013 10112
rect 24228 10084 24501 10112
rect 21968 10072 21974 10084
rect 24489 10081 24501 10084
rect 24535 10112 24547 10115
rect 25498 10112 25504 10124
rect 24535 10084 25504 10112
rect 24535 10081 24547 10084
rect 24489 10075 24547 10081
rect 25498 10072 25504 10084
rect 25556 10072 25562 10124
rect 22462 10044 22468 10056
rect 21836 10016 22468 10044
rect 22462 10004 22468 10016
rect 22520 10004 22526 10056
rect 22649 10047 22707 10053
rect 22649 10013 22661 10047
rect 22695 10044 22707 10047
rect 23474 10044 23480 10056
rect 22695 10016 23480 10044
rect 22695 10013 22707 10016
rect 22649 10007 22707 10013
rect 23474 10004 23480 10016
rect 23532 10004 23538 10056
rect 23750 10004 23756 10056
rect 23808 10044 23814 10056
rect 24765 10047 24823 10053
rect 24765 10044 24777 10047
rect 23808 10016 24777 10044
rect 23808 10004 23814 10016
rect 24765 10013 24777 10016
rect 24811 10013 24823 10047
rect 24765 10007 24823 10013
rect 25774 10004 25780 10056
rect 25832 10044 25838 10056
rect 26973 10047 27031 10053
rect 26973 10044 26985 10047
rect 25832 10016 26985 10044
rect 25832 10004 25838 10016
rect 26973 10013 26985 10016
rect 27019 10013 27031 10047
rect 27430 10044 27436 10056
rect 27391 10016 27436 10044
rect 26973 10007 27031 10013
rect 27430 10004 27436 10016
rect 27488 10004 27494 10056
rect 17586 9936 17592 9988
rect 17644 9976 17650 9988
rect 18141 9979 18199 9985
rect 18141 9976 18153 9979
rect 17644 9948 18153 9976
rect 17644 9936 17650 9948
rect 18141 9945 18153 9948
rect 18187 9945 18199 9979
rect 20042 9979 20100 9985
rect 20042 9976 20054 9979
rect 18141 9939 18199 9945
rect 19536 9948 20054 9976
rect 15528 9880 15884 9908
rect 16025 9911 16083 9917
rect 15528 9868 15534 9880
rect 16025 9877 16037 9911
rect 16071 9908 16083 9911
rect 16574 9908 16580 9920
rect 16071 9880 16580 9908
rect 16071 9877 16083 9880
rect 16025 9871 16083 9877
rect 16574 9868 16580 9880
rect 16632 9868 16638 9920
rect 17865 9911 17923 9917
rect 17865 9877 17877 9911
rect 17911 9908 17923 9911
rect 17954 9908 17960 9920
rect 17911 9880 17960 9908
rect 17911 9877 17923 9880
rect 17865 9871 17923 9877
rect 17954 9868 17960 9880
rect 18012 9868 18018 9920
rect 19536 9917 19564 9948
rect 20042 9945 20054 9948
rect 20088 9945 20100 9979
rect 22916 9979 22974 9985
rect 20042 9939 20100 9945
rect 21192 9948 22876 9976
rect 21192 9920 21220 9948
rect 19521 9911 19579 9917
rect 19521 9877 19533 9911
rect 19567 9877 19579 9911
rect 21174 9908 21180 9920
rect 21135 9880 21180 9908
rect 19521 9871 19579 9877
rect 21174 9868 21180 9880
rect 21232 9868 21238 9920
rect 22002 9908 22008 9920
rect 21963 9880 22008 9908
rect 22002 9868 22008 9880
rect 22060 9868 22066 9920
rect 22848 9908 22876 9948
rect 22916 9945 22928 9979
rect 22962 9976 22974 9979
rect 23014 9976 23020 9988
rect 22962 9948 23020 9976
rect 22962 9945 22974 9948
rect 22916 9939 22974 9945
rect 23014 9936 23020 9948
rect 23072 9936 23078 9988
rect 24486 9976 24492 9988
rect 23860 9948 24492 9976
rect 23860 9908 23888 9948
rect 24486 9936 24492 9948
rect 24544 9936 24550 9988
rect 26728 9979 26786 9985
rect 26728 9945 26740 9979
rect 26774 9976 26786 9979
rect 26774 9948 27292 9976
rect 26774 9945 26786 9948
rect 26728 9939 26786 9945
rect 24026 9908 24032 9920
rect 22848 9880 23888 9908
rect 23939 9880 24032 9908
rect 24026 9868 24032 9880
rect 24084 9908 24090 9920
rect 24673 9911 24731 9917
rect 24673 9908 24685 9911
rect 24084 9880 24685 9908
rect 24084 9868 24090 9880
rect 24673 9877 24685 9880
rect 24719 9877 24731 9911
rect 25130 9908 25136 9920
rect 25091 9880 25136 9908
rect 24673 9871 24731 9877
rect 25130 9868 25136 9880
rect 25188 9868 25194 9920
rect 27264 9917 27292 9948
rect 27249 9911 27307 9917
rect 27249 9877 27261 9911
rect 27295 9877 27307 9911
rect 27249 9871 27307 9877
rect 1104 9818 28888 9840
rect 1104 9766 10214 9818
rect 10266 9766 10278 9818
rect 10330 9766 10342 9818
rect 10394 9766 10406 9818
rect 10458 9766 10470 9818
rect 10522 9766 19478 9818
rect 19530 9766 19542 9818
rect 19594 9766 19606 9818
rect 19658 9766 19670 9818
rect 19722 9766 19734 9818
rect 19786 9766 28888 9818
rect 1104 9744 28888 9766
rect 8507 9707 8565 9713
rect 8507 9704 8519 9707
rect 8220 9676 8519 9704
rect 7742 9636 7748 9648
rect 7208 9608 7748 9636
rect 7208 9577 7236 9608
rect 7742 9596 7748 9608
rect 7800 9596 7806 9648
rect 7929 9639 7987 9645
rect 7929 9605 7941 9639
rect 7975 9636 7987 9639
rect 8220 9636 8248 9676
rect 8507 9673 8519 9676
rect 8553 9704 8565 9707
rect 9122 9704 9128 9716
rect 8553 9676 9128 9704
rect 8553 9673 8565 9676
rect 8507 9667 8565 9673
rect 9122 9664 9128 9676
rect 9180 9664 9186 9716
rect 14734 9704 14740 9716
rect 14695 9676 14740 9704
rect 14734 9664 14740 9676
rect 14792 9664 14798 9716
rect 16758 9704 16764 9716
rect 16719 9676 16764 9704
rect 16758 9664 16764 9676
rect 16816 9664 16822 9716
rect 19889 9707 19947 9713
rect 19889 9673 19901 9707
rect 19935 9704 19947 9707
rect 20070 9704 20076 9716
rect 19935 9676 20076 9704
rect 19935 9673 19947 9676
rect 19889 9667 19947 9673
rect 20070 9664 20076 9676
rect 20128 9664 20134 9716
rect 21821 9707 21879 9713
rect 21821 9673 21833 9707
rect 21867 9704 21879 9707
rect 22002 9704 22008 9716
rect 21867 9676 22008 9704
rect 21867 9673 21879 9676
rect 21821 9667 21879 9673
rect 22002 9664 22008 9676
rect 22060 9664 22066 9716
rect 22462 9664 22468 9716
rect 22520 9704 22526 9716
rect 24026 9704 24032 9716
rect 22520 9676 23888 9704
rect 23987 9676 24032 9704
rect 22520 9664 22526 9676
rect 7975 9608 8248 9636
rect 7975 9605 7987 9608
rect 7929 9599 7987 9605
rect 8294 9596 8300 9648
rect 8352 9636 8358 9648
rect 9306 9636 9312 9648
rect 8352 9608 9312 9636
rect 8352 9596 8358 9608
rect 9306 9596 9312 9608
rect 9364 9596 9370 9648
rect 11146 9596 11152 9648
rect 11204 9636 11210 9648
rect 11885 9639 11943 9645
rect 11885 9636 11897 9639
rect 11204 9608 11897 9636
rect 11204 9596 11210 9608
rect 11885 9605 11897 9608
rect 11931 9605 11943 9639
rect 11885 9599 11943 9605
rect 12253 9639 12311 9645
rect 12253 9605 12265 9639
rect 12299 9636 12311 9639
rect 13078 9636 13084 9648
rect 12299 9608 13084 9636
rect 12299 9605 12311 9608
rect 12253 9599 12311 9605
rect 13078 9596 13084 9608
rect 13136 9596 13142 9648
rect 16209 9639 16267 9645
rect 16209 9605 16221 9639
rect 16255 9636 16267 9639
rect 17678 9636 17684 9648
rect 16255 9608 17684 9636
rect 16255 9605 16267 9608
rect 16209 9599 16267 9605
rect 17678 9596 17684 9608
rect 17736 9596 17742 9648
rect 18138 9596 18144 9648
rect 18196 9636 18202 9648
rect 18294 9639 18352 9645
rect 18294 9636 18306 9639
rect 18196 9608 18306 9636
rect 18196 9596 18202 9608
rect 18294 9605 18306 9608
rect 18340 9605 18352 9639
rect 18294 9599 18352 9605
rect 20349 9639 20407 9645
rect 20349 9605 20361 9639
rect 20395 9636 20407 9639
rect 21174 9636 21180 9648
rect 20395 9608 21180 9636
rect 20395 9605 20407 9608
rect 20349 9599 20407 9605
rect 21174 9596 21180 9608
rect 21232 9596 21238 9648
rect 21453 9639 21511 9645
rect 21453 9605 21465 9639
rect 21499 9636 21511 9639
rect 22554 9636 22560 9648
rect 21499 9608 22560 9636
rect 21499 9605 21511 9608
rect 21453 9599 21511 9605
rect 22554 9596 22560 9608
rect 22612 9596 22618 9648
rect 23860 9636 23888 9676
rect 24026 9664 24032 9676
rect 24084 9664 24090 9716
rect 24670 9704 24676 9716
rect 24631 9676 24676 9704
rect 24670 9664 24676 9676
rect 24728 9664 24734 9716
rect 25130 9704 25136 9716
rect 25091 9676 25136 9704
rect 25130 9664 25136 9676
rect 25188 9664 25194 9716
rect 25961 9707 26019 9713
rect 25961 9673 25973 9707
rect 26007 9704 26019 9707
rect 26142 9704 26148 9716
rect 26007 9676 26148 9704
rect 26007 9673 26019 9676
rect 25961 9667 26019 9673
rect 26142 9664 26148 9676
rect 26200 9664 26206 9716
rect 26421 9707 26479 9713
rect 26421 9673 26433 9707
rect 26467 9704 26479 9707
rect 27430 9704 27436 9716
rect 26467 9676 27436 9704
rect 26467 9673 26479 9676
rect 26421 9667 26479 9673
rect 27430 9664 27436 9676
rect 27488 9664 27494 9716
rect 24946 9636 24952 9648
rect 23860 9608 24952 9636
rect 24946 9596 24952 9608
rect 25004 9596 25010 9648
rect 25041 9639 25099 9645
rect 25041 9605 25053 9639
rect 25087 9636 25099 9639
rect 25682 9636 25688 9648
rect 25087 9608 25688 9636
rect 25087 9605 25099 9608
rect 25041 9599 25099 9605
rect 25682 9596 25688 9608
rect 25740 9596 25746 9648
rect 26050 9636 26056 9648
rect 26011 9608 26056 9636
rect 26050 9596 26056 9608
rect 26108 9596 26114 9648
rect 7193 9571 7251 9577
rect 7193 9537 7205 9571
rect 7239 9537 7251 9571
rect 7193 9531 7251 9537
rect 7374 9528 7380 9580
rect 7432 9568 7438 9580
rect 7469 9571 7527 9577
rect 7469 9568 7481 9571
rect 7432 9540 7481 9568
rect 7432 9528 7438 9540
rect 7469 9537 7481 9540
rect 7515 9568 7527 9571
rect 7837 9571 7895 9577
rect 7837 9568 7849 9571
rect 7515 9540 7849 9568
rect 7515 9537 7527 9540
rect 7469 9531 7527 9537
rect 7837 9537 7849 9540
rect 7883 9537 7895 9571
rect 8018 9568 8024 9580
rect 7979 9540 8024 9568
rect 7837 9531 7895 9537
rect 8018 9528 8024 9540
rect 8076 9528 8082 9580
rect 8662 9568 8668 9580
rect 8496 9540 8668 9568
rect 5813 9503 5871 9509
rect 5813 9469 5825 9503
rect 5859 9500 5871 9503
rect 8496 9500 8524 9540
rect 8662 9528 8668 9540
rect 8720 9528 8726 9580
rect 9030 9568 9036 9580
rect 8991 9540 9036 9568
rect 9030 9528 9036 9540
rect 9088 9528 9094 9580
rect 9122 9528 9128 9580
rect 9180 9568 9186 9580
rect 9766 9577 9772 9580
rect 9217 9571 9275 9577
rect 9217 9568 9229 9571
rect 9180 9540 9229 9568
rect 9180 9528 9186 9540
rect 9217 9537 9229 9540
rect 9263 9537 9275 9571
rect 9760 9568 9772 9577
rect 9727 9540 9772 9568
rect 9217 9531 9275 9537
rect 9760 9531 9772 9540
rect 9766 9528 9772 9531
rect 9824 9528 9830 9580
rect 12069 9571 12127 9577
rect 12069 9537 12081 9571
rect 12115 9568 12127 9571
rect 12526 9568 12532 9580
rect 12115 9540 12434 9568
rect 12487 9540 12532 9568
rect 12115 9537 12127 9540
rect 12069 9531 12127 9537
rect 5859 9472 8524 9500
rect 5859 9469 5871 9472
rect 5813 9463 5871 9469
rect 8846 9460 8852 9512
rect 8904 9460 8910 9512
rect 8938 9460 8944 9512
rect 8996 9500 9002 9512
rect 9493 9503 9551 9509
rect 9493 9500 9505 9503
rect 8996 9472 9505 9500
rect 8996 9460 9002 9472
rect 9493 9469 9505 9472
rect 9539 9469 9551 9503
rect 9493 9463 9551 9469
rect 10502 9460 10508 9512
rect 10560 9500 10566 9512
rect 12250 9500 12256 9512
rect 10560 9472 12256 9500
rect 10560 9460 10566 9472
rect 12250 9460 12256 9472
rect 12308 9460 12314 9512
rect 12406 9500 12434 9540
rect 12526 9528 12532 9540
rect 12584 9528 12590 9580
rect 12710 9568 12716 9580
rect 12671 9540 12716 9568
rect 12710 9528 12716 9540
rect 12768 9528 12774 9580
rect 12802 9528 12808 9580
rect 12860 9568 12866 9580
rect 14001 9571 14059 9577
rect 12860 9540 12905 9568
rect 12860 9528 12866 9540
rect 14001 9537 14013 9571
rect 14047 9568 14059 9571
rect 14458 9568 14464 9580
rect 14047 9540 14464 9568
rect 14047 9537 14059 9540
rect 14001 9531 14059 9537
rect 14458 9528 14464 9540
rect 14516 9528 14522 9580
rect 15838 9528 15844 9580
rect 15896 9568 15902 9580
rect 16117 9571 16175 9577
rect 16117 9568 16129 9571
rect 15896 9540 16129 9568
rect 15896 9528 15902 9540
rect 16117 9537 16129 9540
rect 16163 9537 16175 9571
rect 16298 9568 16304 9580
rect 16259 9540 16304 9568
rect 16117 9531 16175 9537
rect 14090 9500 14096 9512
rect 12406 9472 13768 9500
rect 14051 9472 14096 9500
rect 5537 9435 5595 9441
rect 5537 9401 5549 9435
rect 5583 9432 5595 9435
rect 6914 9432 6920 9444
rect 5583 9404 6920 9432
rect 5583 9401 5595 9404
rect 5537 9395 5595 9401
rect 6914 9392 6920 9404
rect 6972 9392 6978 9444
rect 8864 9432 8892 9460
rect 13740 9444 13768 9472
rect 14090 9460 14096 9472
rect 14148 9500 14154 9512
rect 14553 9503 14611 9509
rect 14553 9500 14565 9503
rect 14148 9472 14565 9500
rect 14148 9460 14154 9472
rect 14553 9469 14565 9472
rect 14599 9469 14611 9503
rect 14553 9463 14611 9469
rect 14737 9503 14795 9509
rect 14737 9469 14749 9503
rect 14783 9469 14795 9503
rect 16132 9500 16160 9531
rect 16298 9528 16304 9540
rect 16356 9528 16362 9580
rect 16669 9571 16727 9577
rect 16669 9568 16681 9571
rect 16408 9540 16681 9568
rect 16408 9500 16436 9540
rect 16669 9537 16681 9540
rect 16715 9537 16727 9571
rect 16669 9531 16727 9537
rect 16853 9571 16911 9577
rect 16853 9537 16865 9571
rect 16899 9537 16911 9571
rect 17310 9568 17316 9580
rect 17271 9540 17316 9568
rect 16853 9531 16911 9537
rect 16132 9472 16436 9500
rect 14737 9463 14795 9469
rect 11146 9432 11152 9444
rect 8864 9404 9251 9432
rect 5353 9367 5411 9373
rect 5353 9333 5365 9367
rect 5399 9364 5411 9367
rect 5994 9364 6000 9376
rect 5399 9336 6000 9364
rect 5399 9333 5411 9336
rect 5353 9327 5411 9333
rect 5994 9324 6000 9336
rect 6052 9324 6058 9376
rect 7009 9367 7067 9373
rect 7009 9333 7021 9367
rect 7055 9364 7067 9367
rect 7098 9364 7104 9376
rect 7055 9336 7104 9364
rect 7055 9333 7067 9336
rect 7009 9327 7067 9333
rect 7098 9324 7104 9336
rect 7156 9324 7162 9376
rect 7377 9367 7435 9373
rect 7377 9333 7389 9367
rect 7423 9364 7435 9367
rect 8018 9364 8024 9376
rect 7423 9336 8024 9364
rect 7423 9333 7435 9336
rect 7377 9327 7435 9333
rect 8018 9324 8024 9336
rect 8076 9324 8082 9376
rect 8478 9364 8484 9376
rect 8439 9336 8484 9364
rect 8478 9324 8484 9336
rect 8536 9324 8542 9376
rect 8662 9324 8668 9376
rect 8720 9364 8726 9376
rect 9223 9364 9251 9404
rect 10704 9404 11152 9432
rect 10704 9364 10732 9404
rect 11146 9392 11152 9404
rect 11204 9432 11210 9444
rect 12342 9432 12348 9444
rect 11204 9404 12348 9432
rect 11204 9392 11210 9404
rect 12342 9392 12348 9404
rect 12400 9392 12406 9444
rect 13722 9392 13728 9444
rect 13780 9432 13786 9444
rect 14752 9432 14780 9463
rect 13780 9404 14780 9432
rect 13780 9392 13786 9404
rect 16298 9392 16304 9444
rect 16356 9432 16362 9444
rect 16868 9432 16896 9531
rect 17310 9528 17316 9540
rect 17368 9528 17374 9580
rect 17402 9528 17408 9580
rect 17460 9568 17466 9580
rect 17460 9540 17505 9568
rect 17460 9528 17466 9540
rect 17586 9528 17592 9580
rect 17644 9568 17650 9580
rect 18046 9568 18052 9580
rect 17644 9540 17689 9568
rect 18007 9540 18052 9568
rect 17644 9528 17650 9540
rect 18046 9528 18052 9540
rect 18104 9528 18110 9580
rect 20257 9571 20315 9577
rect 20257 9568 20269 9571
rect 19076 9540 20269 9568
rect 16356 9404 16896 9432
rect 16356 9392 16362 9404
rect 10870 9364 10876 9376
rect 8720 9336 8765 9364
rect 9223 9336 10732 9364
rect 10831 9336 10876 9364
rect 8720 9324 8726 9336
rect 10870 9324 10876 9336
rect 10928 9324 10934 9376
rect 11238 9324 11244 9376
rect 11296 9364 11302 9376
rect 11422 9364 11428 9376
rect 11296 9336 11428 9364
rect 11296 9324 11302 9336
rect 11422 9324 11428 9336
rect 11480 9324 11486 9376
rect 12434 9324 12440 9376
rect 12492 9364 12498 9376
rect 12529 9367 12587 9373
rect 12529 9364 12541 9367
rect 12492 9336 12541 9364
rect 12492 9324 12498 9336
rect 12529 9333 12541 9336
rect 12575 9333 12587 9367
rect 13630 9364 13636 9376
rect 13591 9336 13636 9364
rect 12529 9327 12587 9333
rect 13630 9324 13636 9336
rect 13688 9324 13694 9376
rect 17589 9367 17647 9373
rect 17589 9333 17601 9367
rect 17635 9364 17647 9367
rect 17770 9364 17776 9376
rect 17635 9336 17776 9364
rect 17635 9333 17647 9336
rect 17589 9327 17647 9333
rect 17770 9324 17776 9336
rect 17828 9324 17834 9376
rect 18230 9324 18236 9376
rect 18288 9364 18294 9376
rect 19076 9364 19104 9540
rect 20257 9537 20269 9540
rect 20303 9537 20315 9571
rect 21266 9568 21272 9580
rect 21227 9540 21272 9568
rect 20257 9531 20315 9537
rect 21266 9528 21272 9540
rect 21324 9528 21330 9580
rect 22186 9528 22192 9580
rect 22244 9568 22250 9580
rect 22934 9571 22992 9577
rect 22934 9568 22946 9571
rect 22244 9540 22946 9568
rect 22244 9528 22250 9540
rect 22934 9537 22946 9540
rect 22980 9537 22992 9571
rect 22934 9531 22992 9537
rect 23201 9571 23259 9577
rect 23201 9537 23213 9571
rect 23247 9568 23259 9571
rect 23382 9568 23388 9580
rect 23247 9540 23388 9568
rect 23247 9537 23259 9540
rect 23201 9531 23259 9537
rect 23382 9528 23388 9540
rect 23440 9528 23446 9580
rect 20530 9500 20536 9512
rect 20491 9472 20536 9500
rect 20530 9460 20536 9472
rect 20588 9460 20594 9512
rect 24121 9503 24179 9509
rect 24121 9469 24133 9503
rect 24167 9469 24179 9503
rect 24121 9463 24179 9469
rect 24305 9503 24363 9509
rect 24305 9469 24317 9503
rect 24351 9500 24363 9503
rect 24854 9500 24860 9512
rect 24351 9472 24860 9500
rect 24351 9469 24363 9472
rect 24305 9463 24363 9469
rect 24026 9392 24032 9444
rect 24084 9432 24090 9444
rect 24136 9432 24164 9463
rect 24854 9460 24860 9472
rect 24912 9500 24918 9512
rect 25225 9503 25283 9509
rect 25225 9500 25237 9503
rect 24912 9472 25237 9500
rect 24912 9460 24918 9472
rect 25225 9469 25237 9472
rect 25271 9469 25283 9503
rect 25225 9463 25283 9469
rect 25777 9503 25835 9509
rect 25777 9469 25789 9503
rect 25823 9469 25835 9503
rect 25777 9463 25835 9469
rect 24084 9404 24164 9432
rect 24084 9392 24090 9404
rect 24946 9392 24952 9444
rect 25004 9432 25010 9444
rect 25792 9432 25820 9463
rect 25004 9404 25820 9432
rect 25004 9392 25010 9404
rect 18288 9336 19104 9364
rect 19429 9367 19487 9373
rect 18288 9324 18294 9336
rect 19429 9333 19441 9367
rect 19475 9364 19487 9367
rect 19702 9364 19708 9376
rect 19475 9336 19708 9364
rect 19475 9333 19487 9336
rect 19429 9327 19487 9333
rect 19702 9324 19708 9336
rect 19760 9324 19766 9376
rect 23658 9364 23664 9376
rect 23619 9336 23664 9364
rect 23658 9324 23664 9336
rect 23716 9324 23722 9376
rect 1104 9274 28888 9296
rect 1104 9222 5582 9274
rect 5634 9222 5646 9274
rect 5698 9222 5710 9274
rect 5762 9222 5774 9274
rect 5826 9222 5838 9274
rect 5890 9222 14846 9274
rect 14898 9222 14910 9274
rect 14962 9222 14974 9274
rect 15026 9222 15038 9274
rect 15090 9222 15102 9274
rect 15154 9222 24110 9274
rect 24162 9222 24174 9274
rect 24226 9222 24238 9274
rect 24290 9222 24302 9274
rect 24354 9222 24366 9274
rect 24418 9222 28888 9274
rect 1104 9200 28888 9222
rect 7374 9160 7380 9172
rect 7335 9132 7380 9160
rect 7374 9120 7380 9132
rect 7432 9120 7438 9172
rect 8478 9120 8484 9172
rect 8536 9160 8542 9172
rect 9214 9160 9220 9172
rect 8536 9132 9220 9160
rect 8536 9120 8542 9132
rect 9214 9120 9220 9132
rect 9272 9120 9278 9172
rect 9766 9120 9772 9172
rect 9824 9160 9830 9172
rect 9953 9163 10011 9169
rect 9953 9160 9965 9163
rect 9824 9132 9965 9160
rect 9824 9120 9830 9132
rect 9953 9129 9965 9132
rect 9999 9129 10011 9163
rect 13630 9160 13636 9172
rect 9953 9123 10011 9129
rect 10888 9132 13636 9160
rect 7392 9024 7420 9120
rect 7837 9095 7895 9101
rect 7837 9061 7849 9095
rect 7883 9092 7895 9095
rect 8018 9092 8024 9104
rect 7883 9064 8024 9092
rect 7883 9061 7895 9064
rect 7837 9055 7895 9061
rect 8018 9052 8024 9064
rect 8076 9052 8082 9104
rect 10042 9024 10048 9036
rect 7392 8996 7696 9024
rect 9955 8996 10048 9024
rect 1854 8956 1860 8968
rect 1815 8928 1860 8956
rect 1854 8916 1860 8928
rect 1912 8916 1918 8968
rect 4614 8916 4620 8968
rect 4672 8956 4678 8968
rect 7668 8965 7696 8996
rect 5997 8959 6055 8965
rect 5997 8956 6009 8959
rect 4672 8928 6009 8956
rect 4672 8916 4678 8928
rect 5997 8925 6009 8928
rect 6043 8956 6055 8959
rect 7653 8959 7711 8965
rect 6043 8928 7604 8956
rect 6043 8925 6055 8928
rect 5997 8919 6055 8925
rect 1670 8888 1676 8900
rect 1631 8860 1676 8888
rect 1670 8848 1676 8860
rect 1728 8888 1734 8900
rect 2133 8891 2191 8897
rect 2133 8888 2145 8891
rect 1728 8860 2145 8888
rect 1728 8848 1734 8860
rect 2133 8857 2145 8860
rect 2179 8857 2191 8891
rect 2133 8851 2191 8857
rect 6264 8891 6322 8897
rect 6264 8857 6276 8891
rect 6310 8888 6322 8891
rect 6822 8888 6828 8900
rect 6310 8860 6828 8888
rect 6310 8857 6322 8860
rect 6264 8851 6322 8857
rect 6822 8848 6828 8860
rect 6880 8848 6886 8900
rect 7576 8888 7604 8928
rect 7653 8925 7665 8959
rect 7699 8925 7711 8959
rect 7653 8919 7711 8925
rect 7926 8916 7932 8968
rect 7984 8965 7990 8968
rect 7984 8959 8033 8965
rect 7984 8925 7987 8959
rect 8021 8925 8033 8959
rect 7984 8919 8033 8925
rect 7984 8916 7990 8919
rect 8110 8916 8116 8968
rect 8168 8956 8174 8968
rect 9968 8965 9996 8996
rect 10042 8984 10048 8996
rect 10100 9024 10106 9036
rect 10502 9024 10508 9036
rect 10100 8996 10508 9024
rect 10100 8984 10106 8996
rect 10502 8984 10508 8996
rect 10560 8984 10566 9036
rect 10888 8965 10916 9132
rect 13630 9120 13636 9132
rect 13688 9120 13694 9172
rect 16669 9163 16727 9169
rect 16669 9129 16681 9163
rect 16715 9160 16727 9163
rect 17310 9160 17316 9172
rect 16715 9132 17316 9160
rect 16715 9129 16727 9132
rect 16669 9123 16727 9129
rect 17310 9120 17316 9132
rect 17368 9120 17374 9172
rect 20441 9163 20499 9169
rect 17420 9132 19334 9160
rect 10962 9052 10968 9104
rect 11020 9052 11026 9104
rect 11514 9092 11520 9104
rect 11164 9064 11520 9092
rect 10986 8965 11014 9052
rect 11164 8965 11192 9064
rect 11514 9052 11520 9064
rect 11572 9052 11578 9104
rect 15286 9092 15292 9104
rect 15247 9064 15292 9092
rect 15286 9052 15292 9064
rect 15344 9052 15350 9104
rect 11422 9024 11428 9036
rect 11256 8996 11428 9024
rect 11256 8965 11284 8996
rect 11422 8984 11428 8996
rect 11480 9024 11486 9036
rect 11882 9024 11888 9036
rect 11480 8996 11888 9024
rect 11480 8984 11486 8996
rect 11882 8984 11888 8996
rect 11940 8984 11946 9036
rect 13998 8984 14004 9036
rect 14056 9024 14062 9036
rect 14056 8996 15148 9024
rect 14056 8984 14062 8996
rect 9953 8959 10011 8965
rect 8168 8928 8213 8956
rect 8168 8916 8174 8928
rect 9953 8925 9965 8959
rect 9999 8925 10011 8959
rect 9953 8919 10011 8925
rect 10229 8959 10287 8965
rect 10229 8925 10241 8959
rect 10275 8956 10287 8959
rect 10689 8959 10747 8965
rect 10689 8956 10701 8959
rect 10275 8928 10701 8956
rect 10275 8925 10287 8928
rect 10229 8919 10287 8925
rect 10689 8925 10701 8928
rect 10735 8925 10747 8959
rect 10689 8919 10747 8925
rect 10873 8959 10931 8965
rect 10873 8925 10885 8959
rect 10919 8925 10931 8959
rect 10986 8959 11055 8965
rect 10986 8928 11009 8959
rect 10873 8919 10931 8925
rect 10997 8925 11009 8928
rect 11043 8925 11055 8959
rect 10997 8919 11055 8925
rect 11149 8959 11207 8965
rect 11149 8925 11161 8959
rect 11195 8925 11207 8959
rect 11149 8919 11207 8925
rect 11241 8959 11299 8965
rect 11241 8925 11253 8959
rect 11287 8925 11299 8959
rect 11241 8919 11299 8925
rect 11348 8928 11928 8956
rect 8386 8888 8392 8900
rect 7576 8860 8392 8888
rect 8386 8848 8392 8860
rect 8444 8848 8450 8900
rect 8570 8848 8576 8900
rect 8628 8888 8634 8900
rect 11348 8888 11376 8928
rect 8628 8860 11376 8888
rect 8628 8848 8634 8860
rect 11422 8848 11428 8900
rect 11480 8888 11486 8900
rect 11609 8891 11667 8897
rect 11609 8888 11621 8891
rect 11480 8860 11621 8888
rect 11480 8848 11486 8860
rect 11609 8857 11621 8860
rect 11655 8857 11667 8891
rect 11609 8851 11667 8857
rect 11793 8891 11851 8897
rect 11793 8857 11805 8891
rect 11839 8857 11851 8891
rect 11900 8888 11928 8928
rect 11974 8916 11980 8968
rect 12032 8956 12038 8968
rect 12434 8965 12440 8968
rect 12161 8959 12219 8965
rect 12161 8956 12173 8959
rect 12032 8928 12173 8956
rect 12032 8916 12038 8928
rect 12161 8925 12173 8928
rect 12207 8925 12219 8959
rect 12161 8919 12219 8925
rect 12428 8919 12440 8965
rect 12492 8956 12498 8968
rect 12492 8928 12528 8956
rect 12434 8916 12440 8919
rect 12492 8916 12498 8928
rect 13630 8916 13636 8968
rect 13688 8956 13694 8968
rect 15013 8959 15071 8965
rect 15013 8956 15025 8959
rect 13688 8928 15025 8956
rect 13688 8916 13694 8928
rect 15013 8925 15025 8928
rect 15059 8925 15071 8959
rect 15120 8956 15148 8996
rect 15194 8984 15200 9036
rect 15252 9024 15258 9036
rect 17420 9024 17448 9132
rect 19306 9092 19334 9132
rect 20441 9129 20453 9163
rect 20487 9160 20499 9163
rect 21266 9160 21272 9172
rect 20487 9132 21272 9160
rect 20487 9129 20499 9132
rect 20441 9123 20499 9129
rect 21266 9120 21272 9132
rect 21324 9160 21330 9172
rect 22097 9163 22155 9169
rect 21324 9132 21956 9160
rect 21324 9120 21330 9132
rect 20990 9092 20996 9104
rect 19306 9064 20996 9092
rect 20990 9052 20996 9064
rect 21048 9052 21054 9104
rect 21726 9092 21732 9104
rect 21687 9064 21732 9092
rect 21726 9052 21732 9064
rect 21784 9052 21790 9104
rect 21928 9092 21956 9132
rect 22097 9129 22109 9163
rect 22143 9160 22155 9163
rect 22186 9160 22192 9172
rect 22143 9132 22192 9160
rect 22143 9129 22155 9132
rect 22097 9123 22155 9129
rect 22186 9120 22192 9132
rect 22244 9120 22250 9172
rect 21928 9064 22094 9092
rect 19702 9024 19708 9036
rect 15252 8996 17448 9024
rect 19663 8996 19708 9024
rect 15252 8984 15258 8996
rect 16960 8965 16988 8996
rect 19702 8984 19708 8996
rect 19760 9024 19766 9036
rect 22066 9024 22094 9064
rect 22373 9027 22431 9033
rect 22373 9024 22385 9027
rect 19760 8996 20300 9024
rect 22066 8996 22385 9024
rect 19760 8984 19766 8996
rect 16853 8959 16911 8965
rect 15120 8950 16804 8956
rect 16853 8950 16865 8959
rect 15120 8928 16865 8950
rect 15013 8919 15071 8925
rect 16776 8925 16865 8928
rect 16899 8925 16911 8959
rect 16776 8922 16911 8925
rect 16853 8919 16911 8922
rect 16945 8959 17003 8965
rect 16945 8925 16957 8959
rect 16991 8925 17003 8959
rect 17129 8959 17187 8965
rect 17129 8956 17141 8959
rect 16945 8919 17003 8925
rect 17052 8928 17141 8956
rect 17052 8900 17080 8928
rect 17129 8925 17141 8928
rect 17175 8925 17187 8959
rect 17129 8919 17187 8925
rect 17221 8959 17279 8965
rect 17221 8925 17233 8959
rect 17267 8925 17279 8959
rect 17221 8919 17279 8925
rect 17497 8959 17555 8965
rect 17497 8925 17509 8959
rect 17543 8956 17555 8959
rect 17586 8956 17592 8968
rect 17543 8928 17592 8956
rect 17543 8925 17555 8928
rect 17497 8919 17555 8925
rect 13814 8888 13820 8900
rect 11900 8860 13820 8888
rect 11793 8851 11851 8857
rect 7650 8820 7656 8832
rect 7611 8792 7656 8820
rect 7650 8780 7656 8792
rect 7708 8780 7714 8832
rect 10134 8820 10140 8832
rect 10095 8792 10140 8820
rect 10134 8780 10140 8792
rect 10192 8780 10198 8832
rect 11808 8820 11836 8851
rect 13814 8848 13820 8860
rect 13872 8848 13878 8900
rect 14458 8848 14464 8900
rect 14516 8888 14522 8900
rect 15105 8891 15163 8897
rect 15105 8888 15117 8891
rect 14516 8860 15117 8888
rect 14516 8848 14522 8860
rect 15105 8857 15117 8860
rect 15151 8888 15163 8891
rect 15194 8888 15200 8900
rect 15151 8860 15200 8888
rect 15151 8857 15163 8860
rect 15105 8851 15163 8857
rect 15194 8848 15200 8860
rect 15252 8848 15258 8900
rect 15289 8891 15347 8897
rect 15289 8857 15301 8891
rect 15335 8888 15347 8891
rect 16666 8888 16672 8900
rect 15335 8860 16672 8888
rect 15335 8857 15347 8860
rect 15289 8851 15347 8857
rect 16666 8848 16672 8860
rect 16724 8848 16730 8900
rect 17034 8848 17040 8900
rect 17092 8848 17098 8900
rect 17236 8888 17264 8919
rect 17586 8916 17592 8928
rect 17644 8916 17650 8968
rect 17770 8965 17776 8968
rect 17764 8956 17776 8965
rect 17731 8928 17776 8956
rect 17764 8919 17776 8928
rect 17770 8916 17776 8919
rect 17828 8916 17834 8968
rect 18230 8916 18236 8968
rect 18288 8956 18294 8968
rect 19337 8959 19395 8965
rect 19337 8956 19349 8959
rect 18288 8928 19349 8956
rect 18288 8916 18294 8928
rect 19337 8925 19349 8928
rect 19383 8925 19395 8959
rect 19886 8956 19892 8968
rect 19799 8928 19892 8956
rect 19337 8919 19395 8925
rect 19886 8916 19892 8928
rect 19944 8956 19950 8968
rect 20272 8958 20300 8996
rect 22373 8993 22385 8996
rect 22419 8993 22431 9027
rect 22373 8987 22431 8993
rect 24854 8984 24860 9036
rect 24912 9024 24918 9036
rect 24949 9027 25007 9033
rect 24949 9024 24961 9027
rect 24912 8996 24961 9024
rect 24912 8984 24918 8996
rect 24949 8993 24961 8996
rect 24995 8993 25007 9027
rect 24949 8987 25007 8993
rect 20349 8959 20407 8965
rect 20349 8958 20361 8959
rect 19944 8928 20015 8956
rect 20272 8930 20361 8958
rect 19944 8916 19950 8928
rect 19987 8888 20015 8928
rect 20349 8925 20361 8930
rect 20395 8925 20407 8959
rect 20349 8919 20407 8925
rect 20533 8959 20591 8965
rect 20533 8925 20545 8959
rect 20579 8956 20591 8959
rect 20714 8956 20720 8968
rect 20579 8928 20720 8956
rect 20579 8925 20591 8928
rect 20533 8919 20591 8925
rect 20714 8916 20720 8928
rect 20772 8916 20778 8968
rect 21634 8916 21640 8968
rect 21692 8956 21698 8968
rect 21821 8959 21879 8965
rect 21692 8928 21737 8956
rect 21692 8916 21698 8928
rect 21821 8925 21833 8959
rect 21867 8925 21879 8959
rect 21821 8919 21879 8925
rect 21913 8959 21971 8965
rect 21913 8925 21925 8959
rect 21959 8956 21971 8959
rect 22002 8956 22008 8968
rect 21959 8928 22008 8956
rect 21959 8925 21971 8928
rect 21913 8919 21971 8925
rect 20438 8888 20444 8900
rect 17236 8860 17908 8888
rect 19987 8860 20444 8888
rect 17880 8832 17908 8860
rect 20438 8848 20444 8860
rect 20496 8848 20502 8900
rect 21836 8832 21864 8919
rect 22002 8916 22008 8928
rect 22060 8916 22066 8968
rect 22649 8959 22707 8965
rect 22649 8925 22661 8959
rect 22695 8956 22707 8959
rect 22830 8956 22836 8968
rect 22695 8928 22836 8956
rect 22695 8925 22707 8928
rect 22649 8919 22707 8925
rect 22830 8916 22836 8928
rect 22888 8916 22894 8968
rect 26053 8959 26111 8965
rect 26053 8956 26065 8959
rect 25608 8928 26065 8956
rect 12066 8820 12072 8832
rect 11808 8792 12072 8820
rect 12066 8780 12072 8792
rect 12124 8780 12130 8832
rect 12250 8780 12256 8832
rect 12308 8820 12314 8832
rect 12434 8820 12440 8832
rect 12308 8792 12440 8820
rect 12308 8780 12314 8792
rect 12434 8780 12440 8792
rect 12492 8780 12498 8832
rect 13078 8780 13084 8832
rect 13136 8820 13142 8832
rect 13541 8823 13599 8829
rect 13541 8820 13553 8823
rect 13136 8792 13553 8820
rect 13136 8780 13142 8792
rect 13541 8789 13553 8792
rect 13587 8789 13599 8823
rect 13541 8783 13599 8789
rect 17862 8780 17868 8832
rect 17920 8820 17926 8832
rect 18877 8823 18935 8829
rect 18877 8820 18889 8823
rect 17920 8792 18889 8820
rect 17920 8780 17926 8792
rect 18877 8789 18889 8792
rect 18923 8789 18935 8823
rect 18877 8783 18935 8789
rect 20073 8823 20131 8829
rect 20073 8789 20085 8823
rect 20119 8820 20131 8823
rect 20530 8820 20536 8832
rect 20119 8792 20536 8820
rect 20119 8789 20131 8792
rect 20073 8783 20131 8789
rect 20530 8780 20536 8792
rect 20588 8780 20594 8832
rect 21818 8780 21824 8832
rect 21876 8780 21882 8832
rect 25130 8820 25136 8832
rect 25091 8792 25136 8820
rect 25130 8780 25136 8792
rect 25188 8780 25194 8832
rect 25222 8780 25228 8832
rect 25280 8820 25286 8832
rect 25608 8829 25636 8928
rect 26053 8925 26065 8928
rect 26099 8925 26111 8959
rect 28350 8956 28356 8968
rect 28311 8928 28356 8956
rect 26053 8919 26111 8925
rect 28350 8916 28356 8928
rect 28408 8916 28414 8968
rect 25593 8823 25651 8829
rect 25280 8792 25325 8820
rect 25280 8780 25286 8792
rect 25593 8789 25605 8823
rect 25639 8789 25651 8823
rect 25866 8820 25872 8832
rect 25827 8792 25872 8820
rect 25593 8783 25651 8789
rect 25866 8780 25872 8792
rect 25924 8780 25930 8832
rect 1104 8730 28888 8752
rect 1104 8678 10214 8730
rect 10266 8678 10278 8730
rect 10330 8678 10342 8730
rect 10394 8678 10406 8730
rect 10458 8678 10470 8730
rect 10522 8678 19478 8730
rect 19530 8678 19542 8730
rect 19594 8678 19606 8730
rect 19658 8678 19670 8730
rect 19722 8678 19734 8730
rect 19786 8678 28888 8730
rect 1104 8656 28888 8678
rect 6822 8616 6828 8628
rect 6783 8588 6828 8616
rect 6822 8576 6828 8588
rect 6880 8576 6886 8628
rect 8021 8619 8079 8625
rect 8021 8585 8033 8619
rect 8067 8616 8079 8619
rect 8478 8616 8484 8628
rect 8067 8588 8484 8616
rect 8067 8585 8079 8588
rect 8021 8579 8079 8585
rect 8478 8576 8484 8588
rect 8536 8616 8542 8628
rect 9490 8616 9496 8628
rect 8536 8588 9496 8616
rect 8536 8576 8542 8588
rect 9490 8576 9496 8588
rect 9548 8576 9554 8628
rect 10134 8576 10140 8628
rect 10192 8616 10198 8628
rect 10413 8619 10471 8625
rect 10413 8616 10425 8619
rect 10192 8588 10425 8616
rect 10192 8576 10198 8588
rect 10413 8585 10425 8588
rect 10459 8585 10471 8619
rect 12713 8619 12771 8625
rect 10413 8579 10471 8585
rect 10520 8588 11560 8616
rect 2041 8551 2099 8557
rect 2041 8517 2053 8551
rect 2087 8548 2099 8551
rect 8570 8548 8576 8560
rect 2087 8520 8576 8548
rect 2087 8517 2099 8520
rect 2041 8511 2099 8517
rect 8570 8508 8576 8520
rect 8628 8508 8634 8560
rect 10520 8548 10548 8588
rect 10336 8520 10548 8548
rect 1394 8440 1400 8492
rect 1452 8480 1458 8492
rect 1673 8483 1731 8489
rect 1673 8480 1685 8483
rect 1452 8452 1685 8480
rect 1452 8440 1458 8452
rect 1673 8449 1685 8452
rect 1719 8449 1731 8483
rect 1673 8443 1731 8449
rect 4884 8483 4942 8489
rect 4884 8449 4896 8483
rect 4930 8480 4942 8483
rect 6362 8480 6368 8492
rect 4930 8452 6368 8480
rect 4930 8449 4942 8452
rect 4884 8443 4942 8449
rect 6362 8440 6368 8452
rect 6420 8440 6426 8492
rect 7098 8480 7104 8492
rect 7059 8452 7104 8480
rect 7098 8440 7104 8452
rect 7156 8440 7162 8492
rect 7837 8483 7895 8489
rect 7837 8449 7849 8483
rect 7883 8449 7895 8483
rect 7837 8443 7895 8449
rect 4614 8412 4620 8424
rect 4575 8384 4620 8412
rect 4614 8372 4620 8384
rect 4672 8372 4678 8424
rect 6825 8415 6883 8421
rect 6825 8381 6837 8415
rect 6871 8412 6883 8415
rect 7650 8412 7656 8424
rect 6871 8384 7656 8412
rect 6871 8381 6883 8384
rect 6825 8375 6883 8381
rect 7650 8372 7656 8384
rect 7708 8372 7714 8424
rect 7852 8344 7880 8443
rect 7926 8440 7932 8492
rect 7984 8480 7990 8492
rect 8113 8483 8171 8489
rect 8113 8480 8125 8483
rect 7984 8452 8125 8480
rect 7984 8440 7990 8452
rect 8113 8449 8125 8452
rect 8159 8449 8171 8483
rect 8386 8480 8392 8492
rect 8347 8452 8392 8480
rect 8113 8443 8171 8449
rect 8386 8440 8392 8452
rect 8444 8440 8450 8492
rect 8656 8483 8714 8489
rect 8656 8449 8668 8483
rect 8702 8480 8714 8483
rect 9674 8480 9680 8492
rect 8702 8452 9680 8480
rect 8702 8449 8714 8452
rect 8656 8443 8714 8449
rect 9674 8440 9680 8452
rect 9732 8440 9738 8492
rect 10045 8483 10103 8489
rect 10045 8480 10057 8483
rect 9784 8452 10057 8480
rect 9784 8353 9812 8452
rect 10045 8449 10057 8452
rect 10091 8449 10103 8483
rect 10045 8443 10103 8449
rect 10183 8483 10241 8489
rect 10183 8449 10195 8483
rect 10229 8480 10241 8483
rect 10336 8480 10364 8520
rect 10686 8508 10692 8560
rect 10744 8548 10750 8560
rect 11422 8548 11428 8560
rect 10744 8520 11428 8548
rect 10744 8508 10750 8520
rect 11422 8508 11428 8520
rect 11480 8508 11486 8560
rect 11532 8492 11560 8588
rect 12713 8585 12725 8619
rect 12759 8616 12771 8619
rect 12802 8616 12808 8628
rect 12759 8588 12808 8616
rect 12759 8585 12771 8588
rect 12713 8579 12771 8585
rect 12802 8576 12808 8588
rect 12860 8576 12866 8628
rect 14093 8619 14151 8625
rect 14093 8585 14105 8619
rect 14139 8616 14151 8619
rect 15838 8616 15844 8628
rect 14139 8588 15844 8616
rect 14139 8585 14151 8588
rect 14093 8579 14151 8585
rect 15838 8576 15844 8588
rect 15896 8576 15902 8628
rect 17402 8576 17408 8628
rect 17460 8616 17466 8628
rect 18049 8619 18107 8625
rect 18049 8616 18061 8619
rect 17460 8588 18061 8616
rect 17460 8576 17466 8588
rect 18049 8585 18061 8588
rect 18095 8585 18107 8619
rect 20070 8616 20076 8628
rect 18049 8579 18107 8585
rect 19168 8588 20076 8616
rect 19168 8560 19196 8588
rect 20070 8576 20076 8588
rect 20128 8616 20134 8628
rect 20714 8616 20720 8628
rect 20128 8588 20720 8616
rect 20128 8576 20134 8588
rect 20714 8576 20720 8588
rect 20772 8576 20778 8628
rect 21634 8576 21640 8628
rect 21692 8616 21698 8628
rect 22465 8619 22523 8625
rect 22465 8616 22477 8619
rect 21692 8588 22477 8616
rect 21692 8576 21698 8588
rect 22465 8585 22477 8588
rect 22511 8585 22523 8619
rect 22465 8579 22523 8585
rect 24857 8619 24915 8625
rect 24857 8585 24869 8619
rect 24903 8616 24915 8619
rect 25222 8616 25228 8628
rect 24903 8588 25228 8616
rect 24903 8585 24915 8588
rect 24857 8579 24915 8585
rect 25222 8576 25228 8588
rect 25280 8576 25286 8628
rect 11793 8551 11851 8557
rect 11793 8517 11805 8551
rect 11839 8548 11851 8551
rect 12161 8551 12219 8557
rect 12161 8548 12173 8551
rect 11839 8520 12173 8548
rect 11839 8517 11851 8520
rect 11793 8511 11851 8517
rect 12161 8517 12173 8520
rect 12207 8517 12219 8551
rect 12161 8511 12219 8517
rect 12345 8551 12403 8557
rect 12345 8517 12357 8551
rect 12391 8548 12403 8551
rect 12434 8548 12440 8560
rect 12391 8520 12440 8548
rect 12391 8517 12403 8520
rect 12345 8511 12403 8517
rect 12434 8508 12440 8520
rect 12492 8548 12498 8560
rect 12894 8548 12900 8560
rect 12492 8520 12900 8548
rect 12492 8508 12498 8520
rect 12894 8508 12900 8520
rect 12952 8508 12958 8560
rect 16206 8548 16212 8560
rect 14568 8520 16212 8548
rect 10229 8452 10364 8480
rect 10229 8449 10241 8452
rect 10183 8443 10241 8449
rect 10410 8440 10416 8492
rect 10468 8480 10474 8492
rect 10505 8483 10563 8489
rect 10505 8480 10517 8483
rect 10468 8452 10517 8480
rect 10468 8440 10474 8452
rect 10505 8449 10517 8452
rect 10551 8449 10563 8483
rect 10505 8443 10563 8449
rect 10594 8440 10600 8492
rect 10652 8480 10658 8492
rect 10781 8483 10839 8489
rect 10781 8480 10793 8483
rect 10652 8452 10793 8480
rect 10652 8440 10658 8452
rect 10781 8449 10793 8452
rect 10827 8449 10839 8483
rect 10781 8443 10839 8449
rect 10870 8440 10876 8492
rect 10928 8480 10934 8492
rect 11514 8480 11520 8492
rect 10928 8452 10973 8480
rect 11475 8452 11520 8480
rect 10928 8440 10934 8452
rect 11514 8440 11520 8452
rect 11572 8440 11578 8492
rect 12066 8480 12072 8492
rect 12027 8452 12072 8480
rect 12066 8440 12072 8452
rect 12124 8440 12130 8492
rect 13078 8480 13084 8492
rect 13039 8452 13084 8480
rect 13078 8440 13084 8452
rect 13136 8440 13142 8492
rect 13262 8480 13268 8492
rect 13223 8452 13268 8480
rect 13262 8440 13268 8452
rect 13320 8440 13326 8492
rect 13449 8483 13507 8489
rect 13449 8449 13461 8483
rect 13495 8480 13507 8483
rect 13998 8480 14004 8492
rect 13495 8452 14004 8480
rect 13495 8449 13507 8452
rect 13449 8443 13507 8449
rect 13998 8440 14004 8452
rect 14056 8440 14062 8492
rect 14274 8480 14280 8492
rect 14235 8452 14280 8480
rect 14274 8440 14280 8452
rect 14332 8440 14338 8492
rect 14458 8480 14464 8492
rect 14419 8452 14464 8480
rect 14458 8440 14464 8452
rect 14516 8440 14522 8492
rect 14568 8489 14596 8520
rect 16206 8508 16212 8520
rect 16264 8508 16270 8560
rect 17034 8508 17040 8560
rect 17092 8548 17098 8560
rect 17681 8551 17739 8557
rect 17681 8548 17693 8551
rect 17092 8520 17693 8548
rect 17092 8508 17098 8520
rect 17681 8517 17693 8520
rect 17727 8517 17739 8551
rect 17681 8511 17739 8517
rect 15194 8489 15200 8492
rect 14553 8483 14611 8489
rect 14553 8449 14565 8483
rect 14599 8449 14611 8483
rect 14553 8443 14611 8449
rect 15188 8443 15200 8489
rect 15252 8480 15258 8492
rect 16224 8480 16252 8508
rect 16853 8483 16911 8489
rect 16853 8480 16865 8483
rect 15252 8452 15288 8480
rect 16224 8452 16865 8480
rect 15194 8440 15200 8443
rect 15252 8440 15258 8452
rect 16853 8449 16865 8452
rect 16899 8480 16911 8483
rect 17313 8483 17371 8489
rect 17313 8480 17325 8483
rect 16899 8452 17325 8480
rect 16899 8449 16911 8452
rect 16853 8443 16911 8449
rect 17313 8449 17325 8452
rect 17359 8449 17371 8483
rect 17313 8443 17371 8449
rect 17497 8483 17555 8489
rect 17497 8449 17509 8483
rect 17543 8449 17555 8483
rect 17696 8480 17724 8511
rect 17862 8508 17868 8560
rect 17920 8548 17926 8560
rect 19150 8548 19156 8560
rect 17920 8520 18184 8548
rect 19063 8520 19156 8548
rect 17920 8508 17926 8520
rect 18156 8489 18184 8520
rect 19150 8508 19156 8520
rect 19208 8508 19214 8560
rect 19337 8551 19395 8557
rect 19337 8517 19349 8551
rect 19383 8548 19395 8551
rect 19426 8548 19432 8560
rect 19383 8520 19432 8548
rect 19383 8517 19395 8520
rect 19337 8511 19395 8517
rect 19426 8508 19432 8520
rect 19484 8548 19490 8560
rect 19886 8548 19892 8560
rect 19484 8520 19892 8548
rect 19484 8508 19490 8520
rect 19886 8508 19892 8520
rect 19944 8508 19950 8560
rect 22646 8548 22652 8560
rect 22607 8520 22652 8548
rect 22646 8508 22652 8520
rect 22704 8508 22710 8560
rect 22830 8548 22836 8560
rect 22791 8520 22836 8548
rect 22830 8508 22836 8520
rect 22888 8508 22894 8560
rect 25492 8551 25550 8557
rect 23492 8520 25268 8548
rect 19978 8489 19984 8492
rect 17957 8483 18015 8489
rect 17957 8480 17969 8483
rect 17696 8452 17969 8480
rect 17497 8443 17555 8449
rect 17957 8449 17969 8452
rect 18003 8449 18015 8483
rect 17957 8443 18015 8449
rect 18141 8483 18199 8489
rect 18141 8449 18153 8483
rect 18187 8449 18199 8483
rect 18141 8443 18199 8449
rect 19972 8443 19984 8489
rect 20036 8480 20042 8492
rect 20036 8452 20072 8480
rect 10321 8415 10379 8421
rect 10321 8381 10333 8415
rect 10367 8412 10379 8415
rect 10686 8412 10692 8424
rect 10367 8384 10692 8412
rect 10367 8381 10379 8384
rect 10321 8375 10379 8381
rect 10686 8372 10692 8384
rect 10744 8372 10750 8424
rect 11790 8412 11796 8424
rect 10796 8384 11796 8412
rect 9769 8347 9827 8353
rect 7852 8316 8432 8344
rect 5997 8279 6055 8285
rect 5997 8245 6009 8279
rect 6043 8276 6055 8279
rect 6086 8276 6092 8288
rect 6043 8248 6092 8276
rect 6043 8245 6055 8248
rect 5997 8239 6055 8245
rect 6086 8236 6092 8248
rect 6144 8236 6150 8288
rect 6914 8236 6920 8288
rect 6972 8276 6978 8288
rect 7009 8279 7067 8285
rect 7009 8276 7021 8279
rect 6972 8248 7021 8276
rect 6972 8236 6978 8248
rect 7009 8245 7021 8248
rect 7055 8276 7067 8279
rect 7650 8276 7656 8288
rect 7055 8248 7656 8276
rect 7055 8245 7067 8248
rect 7009 8239 7067 8245
rect 7650 8236 7656 8248
rect 7708 8236 7714 8288
rect 8404 8276 8432 8316
rect 9769 8313 9781 8347
rect 9815 8344 9827 8347
rect 10502 8344 10508 8356
rect 9815 8316 10508 8344
rect 9815 8313 9827 8316
rect 9769 8307 9827 8313
rect 10502 8304 10508 8316
rect 10560 8344 10566 8356
rect 10796 8344 10824 8384
rect 11790 8372 11796 8384
rect 11848 8372 11854 8424
rect 11882 8372 11888 8424
rect 11940 8412 11946 8424
rect 12250 8412 12256 8424
rect 11940 8384 12256 8412
rect 11940 8372 11946 8384
rect 12250 8372 12256 8384
rect 12308 8412 12314 8424
rect 12989 8415 13047 8421
rect 12989 8412 13001 8415
rect 12308 8384 13001 8412
rect 12308 8372 12314 8384
rect 12989 8381 13001 8384
rect 13035 8381 13047 8415
rect 12989 8375 13047 8381
rect 14090 8372 14096 8424
rect 14148 8412 14154 8424
rect 14369 8415 14427 8421
rect 14369 8412 14381 8415
rect 14148 8384 14381 8412
rect 14148 8372 14154 8384
rect 14369 8381 14381 8384
rect 14415 8381 14427 8415
rect 14369 8375 14427 8381
rect 14734 8372 14740 8424
rect 14792 8412 14798 8424
rect 14921 8415 14979 8421
rect 14921 8412 14933 8415
rect 14792 8384 14933 8412
rect 14792 8372 14798 8384
rect 14921 8381 14933 8384
rect 14967 8381 14979 8415
rect 14921 8375 14979 8381
rect 17037 8415 17095 8421
rect 17037 8381 17049 8415
rect 17083 8412 17095 8415
rect 17512 8412 17540 8443
rect 19978 8440 19984 8443
rect 20036 8440 20042 8452
rect 23492 8424 23520 8520
rect 23750 8489 23756 8492
rect 23744 8443 23756 8489
rect 23808 8480 23814 8492
rect 25240 8489 25268 8520
rect 25492 8517 25504 8551
rect 25538 8548 25550 8551
rect 25866 8548 25872 8560
rect 25538 8520 25872 8548
rect 25538 8517 25550 8520
rect 25492 8511 25550 8517
rect 25866 8508 25872 8520
rect 25924 8508 25930 8560
rect 25225 8483 25283 8489
rect 23808 8452 23844 8480
rect 23750 8440 23756 8443
rect 23808 8440 23814 8452
rect 25225 8449 25237 8483
rect 25271 8449 25283 8483
rect 25225 8443 25283 8449
rect 17083 8384 17540 8412
rect 17083 8381 17095 8384
rect 17037 8375 17095 8381
rect 12342 8344 12348 8356
rect 10560 8316 10824 8344
rect 12303 8316 12348 8344
rect 10560 8304 10566 8316
rect 10686 8276 10692 8288
rect 8404 8248 10692 8276
rect 10686 8236 10692 8248
rect 10744 8236 10750 8288
rect 10796 8285 10824 8316
rect 12342 8304 12348 8316
rect 12400 8304 12406 8356
rect 16301 8347 16359 8353
rect 16301 8313 16313 8347
rect 16347 8344 16359 8347
rect 16942 8344 16948 8356
rect 16347 8316 16948 8344
rect 16347 8313 16359 8316
rect 16301 8307 16359 8313
rect 16942 8304 16948 8316
rect 17000 8344 17006 8356
rect 17052 8344 17080 8375
rect 17586 8372 17592 8424
rect 17644 8412 17650 8424
rect 19705 8415 19763 8421
rect 19705 8412 19717 8415
rect 17644 8384 19717 8412
rect 17644 8372 17650 8384
rect 19705 8381 19717 8384
rect 19751 8381 19763 8415
rect 23474 8412 23480 8424
rect 23435 8384 23480 8412
rect 19705 8375 19763 8381
rect 18690 8344 18696 8356
rect 17000 8316 17080 8344
rect 18651 8316 18696 8344
rect 17000 8304 17006 8316
rect 18690 8304 18696 8316
rect 18748 8344 18754 8356
rect 19334 8344 19340 8356
rect 18748 8316 19340 8344
rect 18748 8304 18754 8316
rect 19334 8304 19340 8316
rect 19392 8304 19398 8356
rect 10781 8279 10839 8285
rect 10781 8245 10793 8279
rect 10827 8245 10839 8279
rect 10781 8239 10839 8245
rect 11149 8279 11207 8285
rect 11149 8245 11161 8279
rect 11195 8276 11207 8279
rect 11238 8276 11244 8288
rect 11195 8248 11244 8276
rect 11195 8245 11207 8248
rect 11149 8239 11207 8245
rect 11238 8236 11244 8248
rect 11296 8236 11302 8288
rect 11606 8276 11612 8288
rect 11567 8248 11612 8276
rect 11606 8236 11612 8248
rect 11664 8236 11670 8288
rect 13170 8276 13176 8288
rect 13131 8248 13176 8276
rect 13170 8236 13176 8248
rect 13228 8236 13234 8288
rect 14182 8236 14188 8288
rect 14240 8276 14246 8288
rect 14458 8276 14464 8288
rect 14240 8248 14464 8276
rect 14240 8236 14246 8248
rect 14458 8236 14464 8248
rect 14516 8236 14522 8288
rect 15562 8236 15568 8288
rect 15620 8276 15626 8288
rect 16669 8279 16727 8285
rect 16669 8276 16681 8279
rect 15620 8248 16681 8276
rect 15620 8236 15626 8248
rect 16669 8245 16681 8248
rect 16715 8245 16727 8279
rect 19720 8276 19748 8375
rect 23474 8372 23480 8384
rect 23532 8372 23538 8424
rect 21082 8344 21088 8356
rect 21043 8316 21088 8344
rect 21082 8304 21088 8316
rect 21140 8304 21146 8356
rect 26605 8347 26663 8353
rect 26605 8344 26617 8347
rect 26160 8316 26617 8344
rect 26160 8288 26188 8316
rect 26605 8313 26617 8316
rect 26651 8313 26663 8347
rect 26605 8307 26663 8313
rect 19886 8276 19892 8288
rect 19720 8248 19892 8276
rect 16669 8239 16727 8245
rect 19886 8236 19892 8248
rect 19944 8236 19950 8288
rect 26142 8236 26148 8288
rect 26200 8236 26206 8288
rect 1104 8186 28888 8208
rect 1104 8134 5582 8186
rect 5634 8134 5646 8186
rect 5698 8134 5710 8186
rect 5762 8134 5774 8186
rect 5826 8134 5838 8186
rect 5890 8134 14846 8186
rect 14898 8134 14910 8186
rect 14962 8134 14974 8186
rect 15026 8134 15038 8186
rect 15090 8134 15102 8186
rect 15154 8134 24110 8186
rect 24162 8134 24174 8186
rect 24226 8134 24238 8186
rect 24290 8134 24302 8186
rect 24354 8134 24366 8186
rect 24418 8134 28888 8186
rect 1104 8112 28888 8134
rect 1394 8072 1400 8084
rect 1355 8044 1400 8072
rect 1394 8032 1400 8044
rect 1452 8032 1458 8084
rect 6362 8072 6368 8084
rect 6323 8044 6368 8072
rect 6362 8032 6368 8044
rect 6420 8032 6426 8084
rect 10410 8032 10416 8084
rect 10468 8072 10474 8084
rect 10689 8075 10747 8081
rect 10689 8072 10701 8075
rect 10468 8044 10701 8072
rect 10468 8032 10474 8044
rect 10689 8041 10701 8044
rect 10735 8072 10747 8075
rect 10870 8072 10876 8084
rect 10735 8044 10876 8072
rect 10735 8041 10747 8044
rect 10689 8035 10747 8041
rect 10870 8032 10876 8044
rect 10928 8032 10934 8084
rect 11514 8072 11520 8084
rect 11475 8044 11520 8072
rect 11514 8032 11520 8044
rect 11572 8032 11578 8084
rect 11977 8075 12035 8081
rect 11977 8041 11989 8075
rect 12023 8072 12035 8075
rect 12066 8072 12072 8084
rect 12023 8044 12072 8072
rect 12023 8041 12035 8044
rect 11977 8035 12035 8041
rect 12066 8032 12072 8044
rect 12124 8032 12130 8084
rect 12437 8075 12495 8081
rect 12437 8041 12449 8075
rect 12483 8072 12495 8075
rect 12710 8072 12716 8084
rect 12483 8044 12716 8072
rect 12483 8041 12495 8044
rect 12437 8035 12495 8041
rect 12710 8032 12716 8044
rect 12768 8032 12774 8084
rect 12894 8032 12900 8084
rect 12952 8072 12958 8084
rect 13265 8075 13323 8081
rect 13265 8072 13277 8075
rect 12952 8044 13277 8072
rect 12952 8032 12958 8044
rect 13265 8041 13277 8044
rect 13311 8041 13323 8075
rect 13265 8035 13323 8041
rect 14182 8032 14188 8084
rect 14240 8072 14246 8084
rect 14277 8075 14335 8081
rect 14277 8072 14289 8075
rect 14240 8044 14289 8072
rect 14240 8032 14246 8044
rect 14277 8041 14289 8044
rect 14323 8041 14335 8075
rect 14277 8035 14335 8041
rect 15105 8075 15163 8081
rect 15105 8041 15117 8075
rect 15151 8072 15163 8075
rect 15194 8072 15200 8084
rect 15151 8044 15200 8072
rect 15151 8041 15163 8044
rect 15105 8035 15163 8041
rect 15194 8032 15200 8044
rect 15252 8032 15258 8084
rect 15286 8032 15292 8084
rect 15344 8072 15350 8084
rect 15473 8075 15531 8081
rect 15473 8072 15485 8075
rect 15344 8044 15485 8072
rect 15344 8032 15350 8044
rect 15473 8041 15485 8044
rect 15519 8041 15531 8075
rect 16206 8072 16212 8084
rect 16167 8044 16212 8072
rect 15473 8035 15531 8041
rect 16206 8032 16212 8044
rect 16264 8032 16270 8084
rect 16482 8072 16488 8084
rect 16443 8044 16488 8072
rect 16482 8032 16488 8044
rect 16540 8032 16546 8084
rect 16942 8072 16948 8084
rect 16903 8044 16948 8072
rect 16942 8032 16948 8044
rect 17000 8032 17006 8084
rect 17957 8075 18015 8081
rect 17957 8041 17969 8075
rect 18003 8072 18015 8075
rect 18046 8072 18052 8084
rect 18003 8044 18052 8072
rect 18003 8041 18015 8044
rect 17957 8035 18015 8041
rect 18046 8032 18052 8044
rect 18104 8072 18110 8084
rect 18322 8072 18328 8084
rect 18104 8044 18328 8072
rect 18104 8032 18110 8044
rect 18322 8032 18328 8044
rect 18380 8032 18386 8084
rect 18506 8032 18512 8084
rect 18564 8072 18570 8084
rect 19245 8075 19303 8081
rect 19245 8072 19257 8075
rect 18564 8044 19257 8072
rect 18564 8032 18570 8044
rect 19245 8041 19257 8044
rect 19291 8041 19303 8075
rect 19245 8035 19303 8041
rect 19978 8032 19984 8084
rect 20036 8072 20042 8084
rect 20073 8075 20131 8081
rect 20073 8072 20085 8075
rect 20036 8044 20085 8072
rect 20036 8032 20042 8044
rect 20073 8041 20085 8044
rect 20119 8041 20131 8075
rect 20622 8072 20628 8084
rect 20073 8035 20131 8041
rect 20180 8044 20628 8072
rect 7006 8004 7012 8016
rect 6104 7976 7012 8004
rect 6104 7948 6132 7976
rect 7006 7964 7012 7976
rect 7064 7964 7070 8016
rect 14093 8007 14151 8013
rect 14093 8004 14105 8007
rect 11532 7976 14105 8004
rect 6086 7936 6092 7948
rect 6047 7908 6092 7936
rect 6086 7896 6092 7908
rect 6144 7896 6150 7948
rect 8113 7939 8171 7945
rect 8113 7936 8125 7939
rect 6564 7908 8125 7936
rect 5813 7871 5871 7877
rect 5813 7837 5825 7871
rect 5859 7837 5871 7871
rect 5813 7831 5871 7837
rect 5828 7800 5856 7831
rect 5902 7828 5908 7880
rect 5960 7868 5966 7880
rect 6564 7877 6592 7908
rect 8113 7905 8125 7908
rect 8159 7905 8171 7939
rect 10502 7936 10508 7948
rect 10463 7908 10508 7936
rect 8113 7899 8171 7905
rect 10502 7896 10508 7908
rect 10560 7896 10566 7948
rect 6914 7877 6920 7880
rect 6549 7871 6607 7877
rect 5960 7840 6005 7868
rect 5960 7828 5966 7840
rect 6549 7837 6561 7871
rect 6595 7837 6607 7871
rect 6549 7831 6607 7837
rect 6871 7871 6920 7877
rect 6871 7837 6883 7871
rect 6917 7837 6920 7871
rect 6871 7831 6920 7837
rect 6914 7828 6920 7831
rect 6972 7828 6978 7880
rect 7006 7828 7012 7880
rect 7064 7868 7070 7880
rect 7558 7868 7564 7880
rect 7064 7840 7109 7868
rect 7519 7840 7564 7868
rect 7064 7828 7070 7840
rect 7558 7828 7564 7840
rect 7616 7828 7622 7880
rect 7745 7871 7803 7877
rect 7745 7837 7757 7871
rect 7791 7868 7803 7871
rect 7834 7868 7840 7880
rect 7791 7840 7840 7868
rect 7791 7837 7803 7840
rect 7745 7831 7803 7837
rect 7834 7828 7840 7840
rect 7892 7828 7898 7880
rect 8018 7868 8024 7880
rect 7979 7840 8024 7868
rect 8018 7828 8024 7840
rect 8076 7828 8082 7880
rect 8205 7871 8263 7877
rect 8205 7837 8217 7871
rect 8251 7837 8263 7871
rect 8205 7831 8263 7837
rect 9585 7871 9643 7877
rect 9585 7837 9597 7871
rect 9631 7868 9643 7871
rect 10042 7868 10048 7880
rect 9631 7840 10048 7868
rect 9631 7837 9643 7840
rect 9585 7831 9643 7837
rect 6454 7800 6460 7812
rect 5828 7772 6460 7800
rect 6454 7760 6460 7772
rect 6512 7760 6518 7812
rect 6638 7800 6644 7812
rect 6599 7772 6644 7800
rect 6638 7760 6644 7772
rect 6696 7760 6702 7812
rect 6730 7760 6736 7812
rect 6788 7800 6794 7812
rect 8220 7800 8248 7831
rect 10042 7828 10048 7840
rect 10100 7828 10106 7880
rect 10413 7871 10471 7877
rect 10413 7837 10425 7871
rect 10459 7868 10471 7871
rect 10594 7868 10600 7880
rect 10459 7840 10600 7868
rect 10459 7837 10471 7840
rect 10413 7831 10471 7837
rect 10594 7828 10600 7840
rect 10652 7828 10658 7880
rect 11532 7877 11560 7976
rect 14093 7973 14105 7976
rect 14139 7973 14151 8007
rect 18598 8004 18604 8016
rect 14093 7967 14151 7973
rect 15856 7976 18604 8004
rect 11701 7939 11759 7945
rect 11701 7905 11713 7939
rect 11747 7936 11759 7939
rect 12434 7936 12440 7948
rect 11747 7908 12440 7936
rect 11747 7905 11759 7908
rect 11701 7899 11759 7905
rect 12434 7896 12440 7908
rect 12492 7896 12498 7948
rect 12529 7939 12587 7945
rect 12529 7905 12541 7939
rect 12575 7936 12587 7939
rect 13078 7936 13084 7948
rect 12575 7908 13084 7936
rect 12575 7905 12587 7908
rect 12529 7899 12587 7905
rect 10689 7871 10747 7877
rect 10689 7837 10701 7871
rect 10735 7868 10747 7871
rect 11517 7871 11575 7877
rect 10735 7840 11468 7868
rect 10735 7837 10747 7840
rect 10689 7831 10747 7837
rect 11054 7800 11060 7812
rect 6788 7772 6833 7800
rect 7576 7772 8248 7800
rect 10520 7772 11060 7800
rect 6788 7760 6794 7772
rect 6089 7735 6147 7741
rect 6089 7701 6101 7735
rect 6135 7732 6147 7735
rect 7576 7732 7604 7772
rect 6135 7704 7604 7732
rect 7653 7735 7711 7741
rect 6135 7701 6147 7704
rect 6089 7695 6147 7701
rect 7653 7701 7665 7735
rect 7699 7732 7711 7735
rect 7834 7732 7840 7744
rect 7699 7704 7840 7732
rect 7699 7701 7711 7704
rect 7653 7695 7711 7701
rect 7834 7692 7840 7704
rect 7892 7692 7898 7744
rect 9953 7735 10011 7741
rect 9953 7701 9965 7735
rect 9999 7732 10011 7735
rect 10520 7732 10548 7772
rect 11054 7760 11060 7772
rect 11112 7760 11118 7812
rect 9999 7704 10548 7732
rect 9999 7701 10011 7704
rect 9953 7695 10011 7701
rect 10686 7692 10692 7744
rect 10744 7732 10750 7744
rect 10873 7735 10931 7741
rect 10873 7732 10885 7735
rect 10744 7704 10885 7732
rect 10744 7692 10750 7704
rect 10873 7701 10885 7704
rect 10919 7701 10931 7735
rect 11440 7732 11468 7840
rect 11517 7837 11529 7871
rect 11563 7837 11575 7871
rect 11790 7868 11796 7880
rect 11751 7840 11796 7868
rect 11517 7831 11575 7837
rect 11790 7828 11796 7840
rect 11848 7828 11854 7880
rect 12250 7868 12256 7880
rect 12211 7840 12256 7868
rect 12250 7828 12256 7840
rect 12308 7828 12314 7880
rect 12345 7871 12403 7877
rect 12345 7837 12357 7871
rect 12391 7837 12403 7871
rect 12345 7831 12403 7837
rect 11606 7760 11612 7812
rect 11664 7800 11670 7812
rect 12360 7800 12388 7831
rect 11664 7772 12388 7800
rect 11664 7760 11670 7772
rect 12544 7732 12572 7899
rect 13078 7896 13084 7908
rect 13136 7896 13142 7948
rect 13354 7896 13360 7948
rect 13412 7936 13418 7948
rect 15562 7936 15568 7948
rect 13412 7908 15332 7936
rect 15523 7908 15568 7936
rect 13412 7896 13418 7908
rect 13262 7828 13268 7880
rect 13320 7868 13326 7880
rect 15304 7877 15332 7908
rect 15562 7896 15568 7908
rect 15620 7896 15626 7948
rect 15856 7877 15884 7976
rect 18598 7964 18604 7976
rect 18656 8004 18662 8016
rect 19610 8004 19616 8016
rect 18656 7976 19616 8004
rect 18656 7964 18662 7976
rect 19610 7964 19616 7976
rect 19668 7964 19674 8016
rect 19705 8007 19763 8013
rect 19705 7973 19717 8007
rect 19751 8004 19763 8007
rect 20180 8004 20208 8044
rect 20622 8032 20628 8044
rect 20680 8032 20686 8084
rect 21177 8075 21235 8081
rect 21177 8041 21189 8075
rect 21223 8072 21235 8075
rect 22278 8072 22284 8084
rect 21223 8044 22284 8072
rect 21223 8041 21235 8044
rect 21177 8035 21235 8041
rect 22278 8032 22284 8044
rect 22336 8032 22342 8084
rect 23750 8072 23756 8084
rect 23711 8044 23756 8072
rect 23750 8032 23756 8044
rect 23808 8032 23814 8084
rect 25130 8032 25136 8084
rect 25188 8072 25194 8084
rect 25317 8075 25375 8081
rect 25317 8072 25329 8075
rect 25188 8044 25329 8072
rect 25188 8032 25194 8044
rect 25317 8041 25329 8044
rect 25363 8041 25375 8075
rect 25317 8035 25375 8041
rect 19751 7976 20208 8004
rect 19751 7973 19763 7976
rect 19705 7967 19763 7973
rect 20530 7964 20536 8016
rect 20588 8004 20594 8016
rect 21726 8004 21732 8016
rect 20588 7976 21732 8004
rect 20588 7964 20594 7976
rect 21726 7964 21732 7976
rect 21784 7964 21790 8016
rect 19150 7936 19156 7948
rect 16592 7908 19156 7936
rect 16592 7877 16620 7908
rect 19150 7896 19156 7908
rect 19208 7896 19214 7948
rect 19334 7936 19340 7948
rect 19295 7908 19340 7936
rect 19334 7896 19340 7908
rect 19392 7896 19398 7948
rect 25866 7936 25872 7948
rect 19536 7908 21404 7936
rect 25827 7908 25872 7936
rect 15289 7871 15347 7877
rect 13320 7840 14504 7868
rect 13320 7828 13326 7840
rect 13357 7803 13415 7809
rect 13357 7769 13369 7803
rect 13403 7800 13415 7803
rect 13630 7800 13636 7812
rect 13403 7772 13636 7800
rect 13403 7769 13415 7772
rect 13357 7763 13415 7769
rect 13630 7760 13636 7772
rect 13688 7760 13694 7812
rect 14274 7809 14280 7812
rect 14261 7803 14280 7809
rect 14261 7769 14273 7803
rect 14261 7763 14280 7769
rect 14274 7760 14280 7763
rect 14332 7760 14338 7812
rect 14476 7809 14504 7840
rect 15289 7837 15301 7871
rect 15335 7868 15347 7871
rect 15841 7871 15899 7877
rect 15841 7868 15853 7871
rect 15335 7840 15853 7868
rect 15335 7837 15347 7840
rect 15289 7831 15347 7837
rect 15841 7837 15853 7840
rect 15887 7837 15899 7871
rect 15841 7831 15899 7837
rect 16485 7871 16543 7877
rect 16485 7837 16497 7871
rect 16531 7837 16543 7871
rect 16485 7831 16543 7837
rect 16577 7871 16635 7877
rect 16577 7837 16589 7871
rect 16623 7837 16635 7871
rect 17034 7868 17040 7880
rect 16577 7831 16635 7837
rect 16684 7840 17040 7868
rect 14461 7803 14519 7809
rect 14461 7769 14473 7803
rect 14507 7769 14519 7803
rect 16500 7800 16528 7831
rect 16684 7800 16712 7840
rect 17034 7828 17040 7840
rect 17092 7828 17098 7880
rect 17129 7871 17187 7877
rect 17129 7837 17141 7871
rect 17175 7868 17187 7871
rect 17862 7868 17868 7880
rect 17175 7840 17868 7868
rect 17175 7837 17187 7840
rect 17129 7831 17187 7837
rect 17862 7828 17868 7840
rect 17920 7828 17926 7880
rect 18322 7828 18328 7880
rect 18380 7868 18386 7880
rect 19536 7877 19564 7908
rect 18693 7871 18751 7877
rect 18693 7868 18705 7871
rect 18380 7840 18705 7868
rect 18380 7828 18386 7840
rect 18693 7837 18705 7840
rect 18739 7837 18751 7871
rect 18693 7831 18751 7837
rect 19521 7871 19579 7877
rect 19521 7837 19533 7871
rect 19567 7837 19579 7871
rect 19521 7831 19579 7837
rect 19610 7828 19616 7880
rect 19668 7868 19674 7880
rect 19978 7868 19984 7880
rect 19668 7840 19984 7868
rect 19668 7828 19674 7840
rect 19978 7828 19984 7840
rect 20036 7868 20042 7880
rect 20257 7871 20315 7877
rect 20257 7868 20269 7871
rect 20036 7840 20269 7868
rect 20036 7828 20042 7840
rect 20257 7837 20269 7840
rect 20303 7837 20315 7871
rect 20438 7868 20444 7880
rect 20399 7840 20444 7868
rect 20257 7831 20315 7837
rect 20438 7828 20444 7840
rect 20496 7828 20502 7880
rect 20530 7828 20536 7880
rect 20588 7868 20594 7880
rect 20809 7871 20867 7877
rect 20588 7840 20633 7868
rect 20588 7828 20594 7840
rect 20809 7837 20821 7871
rect 20855 7868 20867 7871
rect 20990 7868 20996 7880
rect 20855 7840 20996 7868
rect 20855 7837 20867 7840
rect 20809 7831 20867 7837
rect 20990 7828 20996 7840
rect 21048 7828 21054 7880
rect 21269 7871 21327 7877
rect 21269 7868 21281 7871
rect 21100 7840 21281 7868
rect 16500 7772 16712 7800
rect 16853 7803 16911 7809
rect 14461 7763 14519 7769
rect 16853 7769 16865 7803
rect 16899 7769 16911 7803
rect 16853 7763 16911 7769
rect 19245 7803 19303 7809
rect 19245 7769 19257 7803
rect 19291 7800 19303 7803
rect 20622 7800 20628 7812
rect 19291 7772 20628 7800
rect 19291 7769 19303 7772
rect 19245 7763 19303 7769
rect 11440 7704 12572 7732
rect 10873 7695 10931 7701
rect 16482 7692 16488 7744
rect 16540 7732 16546 7744
rect 16868 7732 16896 7763
rect 20622 7760 20628 7772
rect 20680 7760 20686 7812
rect 21100 7800 21128 7840
rect 21269 7837 21281 7840
rect 21315 7837 21327 7871
rect 21376 7868 21404 7908
rect 25866 7896 25872 7908
rect 25924 7896 25930 7948
rect 23017 7871 23075 7877
rect 21376 7840 22968 7868
rect 21269 7831 21327 7837
rect 22750 7803 22808 7809
rect 22750 7800 22762 7803
rect 20732 7772 21128 7800
rect 21284 7772 22762 7800
rect 17310 7732 17316 7744
rect 16540 7704 16896 7732
rect 17271 7704 17316 7732
rect 16540 7692 16546 7704
rect 17310 7692 17316 7704
rect 17368 7692 17374 7744
rect 18325 7735 18383 7741
rect 18325 7701 18337 7735
rect 18371 7732 18383 7735
rect 18506 7732 18512 7744
rect 18371 7704 18512 7732
rect 18371 7701 18383 7704
rect 18325 7695 18383 7701
rect 18506 7692 18512 7704
rect 18564 7692 18570 7744
rect 18785 7735 18843 7741
rect 18785 7701 18797 7735
rect 18831 7732 18843 7735
rect 20254 7732 20260 7744
rect 18831 7704 20260 7732
rect 18831 7701 18843 7704
rect 18785 7695 18843 7701
rect 20254 7692 20260 7704
rect 20312 7732 20318 7744
rect 20732 7732 20760 7772
rect 20898 7732 20904 7744
rect 20312 7704 20760 7732
rect 20859 7704 20904 7732
rect 20312 7692 20318 7704
rect 20898 7692 20904 7704
rect 20956 7692 20962 7744
rect 20993 7735 21051 7741
rect 20993 7701 21005 7735
rect 21039 7732 21051 7735
rect 21174 7732 21180 7744
rect 21039 7704 21180 7732
rect 21039 7701 21051 7704
rect 20993 7695 21051 7701
rect 21174 7692 21180 7704
rect 21232 7692 21238 7744
rect 21284 7741 21312 7772
rect 22750 7769 22762 7772
rect 22796 7769 22808 7803
rect 22940 7800 22968 7840
rect 23017 7837 23029 7871
rect 23063 7868 23075 7871
rect 23474 7868 23480 7880
rect 23063 7840 23480 7868
rect 23063 7837 23075 7840
rect 23017 7831 23075 7837
rect 23474 7828 23480 7840
rect 23532 7828 23538 7880
rect 23569 7871 23627 7877
rect 23569 7837 23581 7871
rect 23615 7868 23627 7871
rect 23658 7868 23664 7880
rect 23615 7840 23664 7868
rect 23615 7837 23627 7840
rect 23569 7831 23627 7837
rect 23658 7828 23664 7840
rect 23716 7828 23722 7880
rect 23934 7828 23940 7880
rect 23992 7868 23998 7880
rect 24397 7871 24455 7877
rect 24397 7868 24409 7871
rect 23992 7840 24409 7868
rect 23992 7828 23998 7840
rect 24397 7837 24409 7840
rect 24443 7837 24455 7871
rect 24397 7831 24455 7837
rect 25406 7828 25412 7880
rect 25464 7868 25470 7880
rect 25777 7871 25835 7877
rect 25777 7868 25789 7871
rect 25464 7840 25789 7868
rect 25464 7828 25470 7840
rect 25777 7837 25789 7840
rect 25823 7868 25835 7871
rect 26142 7868 26148 7880
rect 25823 7840 26148 7868
rect 25823 7837 25835 7840
rect 25777 7831 25835 7837
rect 26142 7828 26148 7840
rect 26200 7828 26206 7880
rect 27893 7871 27951 7877
rect 27893 7837 27905 7871
rect 27939 7868 27951 7871
rect 28350 7868 28356 7880
rect 27939 7840 28356 7868
rect 27939 7837 27951 7840
rect 27893 7831 27951 7837
rect 28350 7828 28356 7840
rect 28408 7828 28414 7880
rect 22940 7772 28212 7800
rect 22750 7763 22808 7769
rect 21269 7735 21327 7741
rect 21269 7701 21281 7735
rect 21315 7701 21327 7735
rect 21269 7695 21327 7701
rect 21358 7692 21364 7744
rect 21416 7732 21422 7744
rect 21637 7735 21695 7741
rect 21637 7732 21649 7735
rect 21416 7704 21649 7732
rect 21416 7692 21422 7704
rect 21637 7701 21649 7704
rect 21683 7701 21695 7735
rect 21637 7695 21695 7701
rect 22646 7692 22652 7744
rect 22704 7732 22710 7744
rect 24489 7735 24547 7741
rect 24489 7732 24501 7735
rect 22704 7704 24501 7732
rect 22704 7692 22710 7704
rect 24489 7701 24501 7704
rect 24535 7701 24547 7735
rect 24489 7695 24547 7701
rect 25685 7735 25743 7741
rect 25685 7701 25697 7735
rect 25731 7732 25743 7735
rect 25774 7732 25780 7744
rect 25731 7704 25780 7732
rect 25731 7701 25743 7704
rect 25685 7695 25743 7701
rect 25774 7692 25780 7704
rect 25832 7692 25838 7744
rect 28184 7741 28212 7772
rect 28169 7735 28227 7741
rect 28169 7701 28181 7735
rect 28215 7701 28227 7735
rect 28169 7695 28227 7701
rect 1104 7642 28888 7664
rect 1104 7590 10214 7642
rect 10266 7590 10278 7642
rect 10330 7590 10342 7642
rect 10394 7590 10406 7642
rect 10458 7590 10470 7642
rect 10522 7590 19478 7642
rect 19530 7590 19542 7642
rect 19594 7590 19606 7642
rect 19658 7590 19670 7642
rect 19722 7590 19734 7642
rect 19786 7590 28888 7642
rect 1104 7568 28888 7590
rect 7469 7531 7527 7537
rect 7469 7497 7481 7531
rect 7515 7497 7527 7531
rect 7469 7491 7527 7497
rect 4884 7463 4942 7469
rect 4884 7429 4896 7463
rect 4930 7460 4942 7463
rect 7484 7460 7512 7491
rect 8110 7488 8116 7540
rect 8168 7528 8174 7540
rect 8757 7531 8815 7537
rect 8757 7528 8769 7531
rect 8168 7500 8769 7528
rect 8168 7488 8174 7500
rect 8757 7497 8769 7500
rect 8803 7528 8815 7531
rect 10962 7528 10968 7540
rect 8803 7500 10968 7528
rect 8803 7497 8815 7500
rect 8757 7491 8815 7497
rect 10962 7488 10968 7500
rect 11020 7488 11026 7540
rect 11882 7488 11888 7540
rect 11940 7528 11946 7540
rect 14458 7528 14464 7540
rect 11940 7500 14464 7528
rect 11940 7488 11946 7500
rect 14458 7488 14464 7500
rect 14516 7528 14522 7540
rect 17402 7528 17408 7540
rect 14516 7500 14780 7528
rect 17363 7500 17408 7528
rect 14516 7488 14522 7500
rect 7834 7460 7840 7472
rect 4930 7432 7512 7460
rect 7795 7432 7840 7460
rect 4930 7429 4942 7432
rect 4884 7423 4942 7429
rect 7834 7420 7840 7432
rect 7892 7420 7898 7472
rect 9309 7463 9367 7469
rect 9309 7429 9321 7463
rect 9355 7460 9367 7463
rect 11054 7460 11060 7472
rect 9355 7432 11060 7460
rect 9355 7429 9367 7432
rect 9309 7423 9367 7429
rect 11054 7420 11060 7432
rect 11112 7420 11118 7472
rect 13262 7460 13268 7472
rect 11624 7432 13268 7460
rect 4614 7392 4620 7404
rect 4575 7364 4620 7392
rect 4614 7352 4620 7364
rect 4672 7352 4678 7404
rect 6365 7395 6423 7401
rect 6365 7361 6377 7395
rect 6411 7392 6423 7395
rect 7006 7392 7012 7404
rect 6411 7364 7012 7392
rect 6411 7361 6423 7364
rect 6365 7355 6423 7361
rect 5997 7259 6055 7265
rect 5997 7225 6009 7259
rect 6043 7256 6055 7259
rect 6380 7256 6408 7355
rect 7006 7352 7012 7364
rect 7064 7352 7070 7404
rect 7650 7392 7656 7404
rect 7611 7364 7656 7392
rect 7650 7352 7656 7364
rect 7708 7352 7714 7404
rect 7745 7395 7803 7401
rect 7745 7361 7757 7395
rect 7791 7361 7803 7395
rect 7745 7355 7803 7361
rect 8021 7395 8079 7401
rect 8021 7361 8033 7395
rect 8067 7392 8079 7395
rect 8478 7392 8484 7404
rect 8067 7364 8484 7392
rect 8067 7361 8079 7364
rect 8021 7355 8079 7361
rect 6454 7284 6460 7336
rect 6512 7324 6518 7336
rect 6641 7327 6699 7333
rect 6641 7324 6653 7327
rect 6512 7296 6653 7324
rect 6512 7284 6518 7296
rect 6641 7293 6653 7296
rect 6687 7324 6699 7327
rect 7558 7324 7564 7336
rect 6687 7296 7564 7324
rect 6687 7293 6699 7296
rect 6641 7287 6699 7293
rect 7558 7284 7564 7296
rect 7616 7324 7622 7336
rect 7760 7324 7788 7355
rect 8478 7352 8484 7364
rect 8536 7352 8542 7404
rect 8665 7395 8723 7401
rect 8665 7361 8677 7395
rect 8711 7392 8723 7395
rect 9769 7395 9827 7401
rect 8711 7364 9720 7392
rect 8711 7361 8723 7364
rect 8665 7355 8723 7361
rect 7616 7296 7788 7324
rect 7616 7284 7622 7296
rect 9122 7256 9128 7268
rect 6043 7228 6408 7256
rect 9083 7228 9128 7256
rect 6043 7225 6055 7228
rect 5997 7219 6055 7225
rect 9122 7216 9128 7228
rect 9180 7216 9186 7268
rect 9692 7256 9720 7364
rect 9769 7361 9781 7395
rect 9815 7392 9827 7395
rect 9858 7392 9864 7404
rect 9815 7364 9864 7392
rect 9815 7361 9827 7364
rect 9769 7355 9827 7361
rect 9858 7352 9864 7364
rect 9916 7352 9922 7404
rect 9953 7395 10011 7401
rect 9953 7361 9965 7395
rect 9999 7361 10011 7395
rect 9953 7355 10011 7361
rect 10321 7395 10379 7401
rect 10321 7361 10333 7395
rect 10367 7392 10379 7395
rect 10502 7392 10508 7404
rect 10367 7364 10508 7392
rect 10367 7361 10379 7364
rect 10321 7355 10379 7361
rect 9968 7324 9996 7355
rect 10502 7352 10508 7364
rect 10560 7352 10566 7404
rect 10597 7395 10655 7401
rect 10597 7361 10609 7395
rect 10643 7392 10655 7395
rect 11146 7392 11152 7404
rect 10643 7364 11152 7392
rect 10643 7361 10655 7364
rect 10597 7355 10655 7361
rect 10612 7324 10640 7355
rect 11146 7352 11152 7364
rect 11204 7392 11210 7404
rect 11514 7392 11520 7404
rect 11204 7364 11520 7392
rect 11204 7352 11210 7364
rect 11514 7352 11520 7364
rect 11572 7352 11578 7404
rect 9968 7296 10640 7324
rect 10778 7284 10784 7336
rect 10836 7324 10842 7336
rect 11624 7324 11652 7432
rect 13262 7420 13268 7432
rect 13320 7460 13326 7472
rect 14752 7460 14780 7500
rect 17402 7488 17408 7500
rect 17460 7488 17466 7540
rect 17494 7488 17500 7540
rect 17552 7488 17558 7540
rect 20898 7488 20904 7540
rect 20956 7528 20962 7540
rect 20956 7500 21956 7528
rect 20956 7488 20962 7500
rect 15470 7460 15476 7472
rect 13320 7432 13676 7460
rect 14752 7432 14872 7460
rect 13320 7420 13326 7432
rect 11793 7395 11851 7401
rect 11793 7361 11805 7395
rect 11839 7392 11851 7395
rect 12434 7392 12440 7404
rect 11839 7364 12440 7392
rect 11839 7361 11851 7364
rect 11793 7355 11851 7361
rect 12406 7352 12440 7364
rect 12492 7352 12498 7404
rect 12618 7352 12624 7404
rect 12676 7392 12682 7404
rect 13648 7401 13676 7432
rect 13357 7395 13415 7401
rect 13357 7392 13369 7395
rect 12676 7364 13369 7392
rect 12676 7352 12682 7364
rect 13357 7361 13369 7364
rect 13403 7361 13415 7395
rect 13357 7355 13415 7361
rect 13633 7395 13691 7401
rect 13633 7361 13645 7395
rect 13679 7361 13691 7395
rect 13633 7355 13691 7361
rect 14366 7352 14372 7404
rect 14424 7392 14430 7404
rect 14844 7401 14872 7432
rect 15120 7432 15476 7460
rect 15120 7401 15148 7432
rect 15470 7420 15476 7432
rect 15528 7460 15534 7472
rect 16482 7460 16488 7472
rect 15528 7432 16488 7460
rect 15528 7420 15534 7432
rect 16482 7420 16488 7432
rect 16540 7420 16546 7472
rect 17221 7463 17279 7469
rect 17221 7429 17233 7463
rect 17267 7460 17279 7463
rect 17512 7460 17540 7488
rect 17267 7432 17540 7460
rect 17267 7429 17279 7432
rect 17221 7423 17279 7429
rect 14737 7395 14795 7401
rect 14737 7392 14749 7395
rect 14424 7364 14749 7392
rect 14424 7352 14430 7364
rect 14737 7361 14749 7364
rect 14783 7361 14795 7395
rect 14737 7355 14795 7361
rect 14829 7395 14887 7401
rect 14829 7361 14841 7395
rect 14875 7361 14887 7395
rect 14829 7355 14887 7361
rect 15013 7395 15071 7401
rect 15013 7361 15025 7395
rect 15059 7361 15071 7395
rect 15013 7355 15071 7361
rect 15105 7395 15163 7401
rect 15105 7361 15117 7395
rect 15151 7361 15163 7395
rect 15838 7392 15844 7404
rect 15799 7364 15844 7392
rect 15105 7355 15163 7361
rect 10836 7296 11652 7324
rect 10836 7284 10842 7296
rect 12158 7284 12164 7336
rect 12216 7324 12222 7336
rect 12253 7327 12311 7333
rect 12253 7324 12265 7327
rect 12216 7296 12265 7324
rect 12216 7284 12222 7296
rect 12253 7293 12265 7296
rect 12299 7293 12311 7327
rect 12406 7324 12434 7352
rect 12529 7327 12587 7333
rect 12529 7324 12541 7327
rect 12406 7296 12541 7324
rect 12253 7287 12311 7293
rect 12529 7293 12541 7296
rect 12575 7324 12587 7327
rect 13170 7324 13176 7336
rect 12575 7296 13176 7324
rect 12575 7293 12587 7296
rect 12529 7287 12587 7293
rect 9766 7256 9772 7268
rect 9679 7228 9772 7256
rect 9766 7216 9772 7228
rect 9824 7256 9830 7268
rect 10796 7256 10824 7284
rect 9824 7228 10824 7256
rect 12268 7256 12296 7287
rect 13170 7284 13176 7296
rect 13228 7284 13234 7336
rect 14642 7284 14648 7336
rect 14700 7324 14706 7336
rect 15028 7324 15056 7355
rect 15838 7352 15844 7364
rect 15896 7352 15902 7404
rect 15930 7352 15936 7404
rect 15988 7392 15994 7404
rect 16117 7395 16175 7401
rect 15988 7364 16033 7392
rect 15988 7352 15994 7364
rect 16117 7361 16129 7395
rect 16163 7392 16175 7395
rect 17034 7392 17040 7404
rect 16163 7364 17040 7392
rect 16163 7361 16175 7364
rect 16117 7355 16175 7361
rect 17034 7352 17040 7364
rect 17092 7392 17098 7404
rect 17236 7392 17264 7423
rect 19978 7420 19984 7472
rect 20036 7460 20042 7472
rect 20530 7460 20536 7472
rect 20036 7432 20536 7460
rect 20036 7420 20042 7432
rect 20530 7420 20536 7432
rect 20588 7420 20594 7472
rect 20990 7460 20996 7472
rect 20951 7432 20996 7460
rect 20990 7420 20996 7432
rect 21048 7420 21054 7472
rect 21174 7420 21180 7472
rect 21232 7460 21238 7472
rect 21818 7460 21824 7472
rect 21232 7432 21824 7460
rect 21232 7420 21238 7432
rect 21818 7420 21824 7432
rect 21876 7420 21882 7472
rect 21928 7469 21956 7500
rect 24026 7488 24032 7540
rect 24084 7528 24090 7540
rect 24121 7531 24179 7537
rect 24121 7528 24133 7531
rect 24084 7500 24133 7528
rect 24084 7488 24090 7500
rect 24121 7497 24133 7500
rect 24167 7497 24179 7531
rect 24121 7491 24179 7497
rect 24581 7531 24639 7537
rect 24581 7497 24593 7531
rect 24627 7528 24639 7531
rect 25222 7528 25228 7540
rect 24627 7500 25228 7528
rect 24627 7497 24639 7500
rect 24581 7491 24639 7497
rect 25222 7488 25228 7500
rect 25280 7488 25286 7540
rect 21913 7463 21971 7469
rect 21913 7429 21925 7463
rect 21959 7460 21971 7463
rect 22646 7460 22652 7472
rect 21959 7432 22652 7460
rect 21959 7429 21971 7432
rect 21913 7423 21971 7429
rect 22646 7420 22652 7432
rect 22704 7420 22710 7472
rect 22865 7463 22923 7469
rect 22865 7429 22877 7463
rect 22911 7460 22923 7463
rect 24486 7460 24492 7472
rect 22911 7432 23796 7460
rect 24447 7432 24492 7460
rect 22911 7429 22923 7432
rect 22865 7423 22923 7429
rect 17494 7392 17500 7404
rect 17092 7364 17264 7392
rect 17455 7364 17500 7392
rect 17092 7352 17098 7364
rect 17494 7352 17500 7364
rect 17552 7352 17558 7404
rect 17586 7352 17592 7404
rect 17644 7392 17650 7404
rect 17773 7395 17831 7401
rect 17773 7392 17785 7395
rect 17644 7364 17785 7392
rect 17644 7352 17650 7364
rect 17773 7361 17785 7364
rect 17819 7361 17831 7395
rect 18029 7395 18087 7401
rect 18029 7392 18041 7395
rect 17773 7355 17831 7361
rect 17880 7364 18041 7392
rect 17880 7324 17908 7364
rect 18029 7361 18041 7364
rect 18075 7361 18087 7395
rect 18029 7355 18087 7361
rect 19334 7352 19340 7404
rect 19392 7392 19398 7404
rect 19613 7395 19671 7401
rect 19613 7392 19625 7395
rect 19392 7364 19625 7392
rect 19392 7352 19398 7364
rect 19613 7361 19625 7364
rect 19659 7392 19671 7395
rect 19702 7392 19708 7404
rect 19659 7364 19708 7392
rect 19659 7361 19671 7364
rect 19613 7355 19671 7361
rect 19702 7352 19708 7364
rect 19760 7352 19766 7404
rect 20806 7392 20812 7404
rect 20767 7364 20812 7392
rect 20806 7352 20812 7364
rect 20864 7352 20870 7404
rect 23385 7395 23443 7401
rect 23385 7392 23397 7395
rect 22066 7364 23397 7392
rect 14700 7296 15056 7324
rect 17236 7296 17908 7324
rect 19889 7327 19947 7333
rect 14700 7284 14706 7296
rect 12894 7256 12900 7268
rect 12268 7228 12900 7256
rect 9824 7216 9830 7228
rect 12894 7216 12900 7228
rect 12952 7216 12958 7268
rect 17236 7265 17264 7296
rect 19889 7293 19901 7327
rect 19935 7324 19947 7327
rect 19978 7324 19984 7336
rect 19935 7296 19984 7324
rect 19935 7293 19947 7296
rect 19889 7287 19947 7293
rect 19978 7284 19984 7296
rect 20036 7284 20042 7336
rect 21634 7284 21640 7336
rect 21692 7324 21698 7336
rect 22066 7324 22094 7364
rect 23385 7361 23397 7364
rect 23431 7361 23443 7395
rect 23768 7392 23796 7432
rect 24486 7420 24492 7432
rect 24544 7420 24550 7472
rect 24946 7460 24952 7472
rect 24596 7432 24952 7460
rect 24596 7392 24624 7432
rect 24946 7420 24952 7432
rect 25004 7420 25010 7472
rect 23768 7364 24624 7392
rect 23385 7355 23443 7361
rect 24854 7352 24860 7404
rect 24912 7392 24918 7404
rect 25317 7395 25375 7401
rect 25317 7392 25329 7395
rect 24912 7364 25329 7392
rect 24912 7352 24918 7364
rect 25317 7361 25329 7364
rect 25363 7361 25375 7395
rect 25317 7355 25375 7361
rect 21692 7296 22094 7324
rect 22189 7327 22247 7333
rect 21692 7284 21698 7296
rect 22189 7293 22201 7327
rect 22235 7293 22247 7327
rect 22189 7287 22247 7293
rect 17221 7259 17279 7265
rect 17221 7225 17233 7259
rect 17267 7225 17279 7259
rect 17221 7219 17279 7225
rect 21358 7216 21364 7268
rect 21416 7256 21422 7268
rect 22204 7256 22232 7287
rect 22278 7284 22284 7336
rect 22336 7324 22342 7336
rect 22336 7296 22381 7324
rect 22336 7284 22342 7296
rect 22830 7284 22836 7336
rect 22888 7324 22894 7336
rect 24673 7327 24731 7333
rect 24673 7324 24685 7327
rect 22888 7296 24685 7324
rect 22888 7284 22894 7296
rect 24673 7293 24685 7296
rect 24719 7324 24731 7327
rect 25501 7327 25559 7333
rect 25501 7324 25513 7327
rect 24719 7296 25513 7324
rect 24719 7293 24731 7296
rect 24673 7287 24731 7293
rect 25501 7293 25513 7296
rect 25547 7324 25559 7327
rect 25866 7324 25872 7336
rect 25547 7296 25872 7324
rect 25547 7293 25559 7296
rect 25501 7287 25559 7293
rect 25866 7284 25872 7296
rect 25924 7284 25930 7336
rect 23566 7256 23572 7268
rect 21416 7228 22232 7256
rect 23527 7228 23572 7256
rect 21416 7216 21422 7228
rect 23566 7216 23572 7228
rect 23624 7216 23630 7268
rect 9858 7188 9864 7200
rect 9819 7160 9864 7188
rect 9858 7148 9864 7160
rect 9916 7148 9922 7200
rect 9950 7148 9956 7200
rect 10008 7188 10014 7200
rect 11606 7188 11612 7200
rect 10008 7160 11612 7188
rect 10008 7148 10014 7160
rect 11606 7148 11612 7160
rect 11664 7188 11670 7200
rect 11885 7191 11943 7197
rect 11885 7188 11897 7191
rect 11664 7160 11897 7188
rect 11664 7148 11670 7160
rect 11885 7157 11897 7160
rect 11931 7157 11943 7191
rect 11885 7151 11943 7157
rect 14366 7148 14372 7200
rect 14424 7188 14430 7200
rect 14553 7191 14611 7197
rect 14553 7188 14565 7191
rect 14424 7160 14565 7188
rect 14424 7148 14430 7160
rect 14553 7157 14565 7160
rect 14599 7157 14611 7191
rect 14553 7151 14611 7157
rect 16022 7148 16028 7200
rect 16080 7188 16086 7200
rect 16117 7191 16175 7197
rect 16117 7188 16129 7191
rect 16080 7160 16129 7188
rect 16080 7148 16086 7160
rect 16117 7157 16129 7160
rect 16163 7157 16175 7191
rect 16117 7151 16175 7157
rect 18414 7148 18420 7200
rect 18472 7188 18478 7200
rect 19058 7188 19064 7200
rect 18472 7160 19064 7188
rect 18472 7148 18478 7160
rect 19058 7148 19064 7160
rect 19116 7188 19122 7200
rect 19153 7191 19211 7197
rect 19153 7188 19165 7191
rect 19116 7160 19165 7188
rect 19116 7148 19122 7160
rect 19153 7157 19165 7160
rect 19199 7157 19211 7191
rect 19153 7151 19211 7157
rect 21726 7148 21732 7200
rect 21784 7188 21790 7200
rect 22097 7191 22155 7197
rect 22097 7188 22109 7191
rect 21784 7160 22109 7188
rect 21784 7148 21790 7160
rect 22097 7157 22109 7160
rect 22143 7157 22155 7191
rect 22830 7188 22836 7200
rect 22791 7160 22836 7188
rect 22097 7151 22155 7157
rect 22830 7148 22836 7160
rect 22888 7148 22894 7200
rect 23017 7191 23075 7197
rect 23017 7157 23029 7191
rect 23063 7188 23075 7191
rect 23106 7188 23112 7200
rect 23063 7160 23112 7188
rect 23063 7157 23075 7160
rect 23017 7151 23075 7157
rect 23106 7148 23112 7160
rect 23164 7148 23170 7200
rect 25133 7191 25191 7197
rect 25133 7157 25145 7191
rect 25179 7188 25191 7191
rect 25314 7188 25320 7200
rect 25179 7160 25320 7188
rect 25179 7157 25191 7160
rect 25133 7151 25191 7157
rect 25314 7148 25320 7160
rect 25372 7148 25378 7200
rect 1104 7098 28888 7120
rect 1104 7046 5582 7098
rect 5634 7046 5646 7098
rect 5698 7046 5710 7098
rect 5762 7046 5774 7098
rect 5826 7046 5838 7098
rect 5890 7046 14846 7098
rect 14898 7046 14910 7098
rect 14962 7046 14974 7098
rect 15026 7046 15038 7098
rect 15090 7046 15102 7098
rect 15154 7046 24110 7098
rect 24162 7046 24174 7098
rect 24226 7046 24238 7098
rect 24290 7046 24302 7098
rect 24354 7046 24366 7098
rect 24418 7046 28888 7098
rect 1104 7024 28888 7046
rect 5902 6944 5908 6996
rect 5960 6984 5966 6996
rect 6917 6987 6975 6993
rect 6917 6984 6929 6987
rect 5960 6956 6929 6984
rect 5960 6944 5966 6956
rect 6917 6953 6929 6956
rect 6963 6984 6975 6987
rect 7098 6984 7104 6996
rect 6963 6956 7104 6984
rect 6963 6953 6975 6956
rect 6917 6947 6975 6953
rect 7098 6944 7104 6956
rect 7156 6944 7162 6996
rect 7285 6987 7343 6993
rect 7285 6953 7297 6987
rect 7331 6984 7343 6987
rect 8018 6984 8024 6996
rect 7331 6956 8024 6984
rect 7331 6953 7343 6956
rect 7285 6947 7343 6953
rect 8018 6944 8024 6956
rect 8076 6944 8082 6996
rect 8386 6944 8392 6996
rect 8444 6984 8450 6996
rect 8570 6984 8576 6996
rect 8444 6956 8576 6984
rect 8444 6944 8450 6956
rect 8570 6944 8576 6956
rect 8628 6984 8634 6996
rect 9122 6984 9128 6996
rect 8628 6956 9128 6984
rect 8628 6944 8634 6956
rect 4614 6876 4620 6928
rect 4672 6916 4678 6928
rect 4672 6888 5580 6916
rect 4672 6876 4678 6888
rect 5552 6780 5580 6888
rect 7926 6876 7932 6928
rect 7984 6916 7990 6928
rect 7984 6888 8524 6916
rect 7984 6876 7990 6888
rect 6641 6783 6699 6789
rect 6641 6780 6653 6783
rect 5552 6752 6653 6780
rect 6641 6749 6653 6752
rect 6687 6749 6699 6783
rect 6914 6780 6920 6792
rect 6875 6752 6920 6780
rect 6641 6743 6699 6749
rect 6914 6740 6920 6752
rect 6972 6740 6978 6792
rect 7006 6740 7012 6792
rect 7064 6780 7070 6792
rect 7926 6780 7932 6792
rect 7064 6752 7109 6780
rect 7887 6752 7932 6780
rect 7064 6740 7070 6752
rect 7926 6740 7932 6752
rect 7984 6740 7990 6792
rect 8021 6783 8079 6789
rect 8021 6749 8033 6783
rect 8067 6749 8079 6783
rect 8021 6743 8079 6749
rect 8205 6783 8263 6789
rect 8205 6749 8217 6783
rect 8251 6749 8263 6783
rect 8205 6743 8263 6749
rect 8297 6783 8355 6789
rect 8297 6749 8309 6783
rect 8343 6780 8355 6783
rect 8386 6780 8392 6792
rect 8343 6752 8392 6780
rect 8343 6749 8355 6752
rect 8297 6743 8355 6749
rect 6362 6712 6368 6724
rect 6420 6721 6426 6724
rect 6332 6684 6368 6712
rect 6362 6672 6368 6684
rect 6420 6675 6432 6721
rect 6420 6672 6426 6675
rect 5261 6647 5319 6653
rect 5261 6613 5273 6647
rect 5307 6644 5319 6647
rect 5902 6644 5908 6656
rect 5307 6616 5908 6644
rect 5307 6613 5319 6616
rect 5261 6607 5319 6613
rect 5902 6604 5908 6616
rect 5960 6604 5966 6656
rect 7742 6644 7748 6656
rect 7703 6616 7748 6644
rect 7742 6604 7748 6616
rect 7800 6604 7806 6656
rect 8036 6644 8064 6743
rect 8220 6712 8248 6743
rect 8386 6740 8392 6752
rect 8444 6740 8450 6792
rect 8496 6780 8524 6888
rect 8956 6857 8984 6956
rect 9122 6944 9128 6956
rect 9180 6944 9186 6996
rect 9214 6944 9220 6996
rect 9272 6984 9278 6996
rect 10321 6987 10379 6993
rect 9272 6956 9904 6984
rect 9272 6944 9278 6956
rect 9876 6916 9904 6956
rect 10321 6953 10333 6987
rect 10367 6984 10379 6987
rect 10502 6984 10508 6996
rect 10367 6956 10508 6984
rect 10367 6953 10379 6956
rect 10321 6947 10379 6953
rect 10502 6944 10508 6956
rect 10560 6944 10566 6996
rect 12526 6984 12532 6996
rect 10612 6956 12532 6984
rect 10612 6916 10640 6956
rect 12526 6944 12532 6956
rect 12584 6944 12590 6996
rect 15470 6984 15476 6996
rect 15431 6956 15476 6984
rect 15470 6944 15476 6956
rect 15528 6944 15534 6996
rect 17402 6944 17408 6996
rect 17460 6984 17466 6996
rect 17589 6987 17647 6993
rect 17589 6984 17601 6987
rect 17460 6956 17601 6984
rect 17460 6944 17466 6956
rect 17589 6953 17601 6956
rect 17635 6953 17647 6987
rect 18414 6984 18420 6996
rect 18375 6956 18420 6984
rect 17589 6947 17647 6953
rect 18414 6944 18420 6956
rect 18472 6944 18478 6996
rect 20530 6984 20536 6996
rect 20491 6956 20536 6984
rect 20530 6944 20536 6956
rect 20588 6944 20594 6996
rect 23934 6944 23940 6996
rect 23992 6984 23998 6996
rect 24029 6987 24087 6993
rect 24029 6984 24041 6987
rect 23992 6956 24041 6984
rect 23992 6944 23998 6956
rect 24029 6953 24041 6956
rect 24075 6953 24087 6987
rect 24029 6947 24087 6953
rect 12158 6916 12164 6928
rect 9876 6888 10640 6916
rect 12119 6888 12164 6916
rect 12158 6876 12164 6888
rect 12216 6876 12222 6928
rect 12253 6919 12311 6925
rect 12253 6885 12265 6919
rect 12299 6885 12311 6919
rect 12253 6879 12311 6885
rect 8941 6851 8999 6857
rect 8941 6817 8953 6851
rect 8987 6817 8999 6851
rect 11882 6848 11888 6860
rect 8941 6811 8999 6817
rect 10888 6820 11888 6848
rect 10778 6780 10784 6792
rect 8496 6752 9812 6780
rect 10739 6752 10784 6780
rect 9208 6715 9266 6721
rect 8220 6684 9168 6712
rect 8294 6644 8300 6656
rect 8036 6616 8300 6644
rect 8294 6604 8300 6616
rect 8352 6604 8358 6656
rect 9140 6644 9168 6684
rect 9208 6681 9220 6715
rect 9254 6712 9266 6715
rect 9674 6712 9680 6724
rect 9254 6684 9680 6712
rect 9254 6681 9266 6684
rect 9208 6675 9266 6681
rect 9674 6672 9680 6684
rect 9732 6672 9738 6724
rect 9784 6712 9812 6752
rect 10778 6740 10784 6752
rect 10836 6740 10842 6792
rect 10888 6789 10916 6820
rect 11882 6808 11888 6820
rect 11940 6808 11946 6860
rect 12268 6848 12296 6879
rect 17494 6876 17500 6928
rect 17552 6916 17558 6928
rect 17957 6919 18015 6925
rect 17957 6916 17969 6919
rect 17552 6888 17969 6916
rect 17552 6876 17558 6888
rect 17957 6885 17969 6888
rect 18003 6885 18015 6919
rect 17957 6879 18015 6885
rect 11992 6820 12296 6848
rect 10873 6783 10931 6789
rect 10873 6749 10885 6783
rect 10919 6749 10931 6783
rect 10873 6743 10931 6749
rect 11057 6783 11115 6789
rect 11057 6749 11069 6783
rect 11103 6749 11115 6783
rect 11057 6743 11115 6749
rect 11072 6712 11100 6743
rect 11146 6740 11152 6792
rect 11204 6780 11210 6792
rect 11204 6752 11249 6780
rect 11204 6740 11210 6752
rect 11330 6740 11336 6792
rect 11388 6780 11394 6792
rect 11517 6783 11575 6789
rect 11517 6780 11529 6783
rect 11388 6752 11529 6780
rect 11388 6740 11394 6752
rect 11517 6749 11529 6752
rect 11563 6780 11575 6783
rect 11698 6780 11704 6792
rect 11563 6752 11704 6780
rect 11563 6749 11575 6752
rect 11517 6743 11575 6749
rect 11698 6740 11704 6752
rect 11756 6740 11762 6792
rect 11422 6712 11428 6724
rect 9784 6684 10732 6712
rect 11072 6684 11428 6712
rect 10042 6644 10048 6656
rect 9140 6616 10048 6644
rect 10042 6604 10048 6616
rect 10100 6604 10106 6656
rect 10594 6644 10600 6656
rect 10555 6616 10600 6644
rect 10594 6604 10600 6616
rect 10652 6604 10658 6656
rect 10704 6644 10732 6684
rect 11422 6672 11428 6684
rect 11480 6712 11486 6724
rect 11992 6712 12020 6820
rect 17310 6808 17316 6860
rect 17368 6848 17374 6860
rect 17681 6851 17739 6857
rect 17368 6820 17540 6848
rect 17368 6808 17374 6820
rect 12069 6783 12127 6789
rect 12069 6749 12081 6783
rect 12115 6749 12127 6783
rect 12069 6743 12127 6749
rect 12381 6783 12439 6789
rect 12381 6749 12393 6783
rect 12427 6780 12439 6783
rect 12710 6780 12716 6792
rect 12427 6752 12716 6780
rect 12427 6749 12439 6752
rect 12381 6743 12439 6749
rect 11480 6684 12020 6712
rect 11480 6672 11486 6684
rect 11330 6644 11336 6656
rect 10704 6616 11336 6644
rect 11330 6604 11336 6616
rect 11388 6604 11394 6656
rect 11790 6604 11796 6656
rect 11848 6644 11854 6656
rect 11885 6647 11943 6653
rect 11885 6644 11897 6647
rect 11848 6616 11897 6644
rect 11848 6604 11854 6616
rect 11885 6613 11897 6616
rect 11931 6613 11943 6647
rect 12084 6644 12112 6743
rect 12710 6740 12716 6752
rect 12768 6740 12774 6792
rect 12894 6780 12900 6792
rect 12855 6752 12900 6780
rect 12894 6740 12900 6752
rect 12952 6740 12958 6792
rect 13630 6780 13636 6792
rect 13591 6752 13636 6780
rect 13630 6740 13636 6752
rect 13688 6740 13694 6792
rect 13906 6740 13912 6792
rect 13964 6780 13970 6792
rect 14093 6783 14151 6789
rect 14093 6780 14105 6783
rect 13964 6752 14105 6780
rect 13964 6740 13970 6752
rect 14093 6749 14105 6752
rect 14139 6780 14151 6783
rect 14734 6780 14740 6792
rect 14139 6752 14740 6780
rect 14139 6749 14151 6752
rect 14093 6743 14151 6749
rect 14734 6740 14740 6752
rect 14792 6780 14798 6792
rect 16022 6789 16028 6792
rect 15749 6783 15807 6789
rect 15749 6780 15761 6783
rect 14792 6752 15761 6780
rect 14792 6740 14798 6752
rect 15749 6749 15761 6752
rect 15795 6749 15807 6783
rect 16016 6780 16028 6789
rect 15983 6752 16028 6780
rect 15749 6743 15807 6749
rect 16016 6743 16028 6752
rect 16022 6740 16028 6743
rect 16080 6740 16086 6792
rect 17512 6789 17540 6820
rect 17681 6817 17693 6851
rect 17727 6848 17739 6851
rect 18432 6848 18460 6944
rect 20073 6919 20131 6925
rect 20073 6885 20085 6919
rect 20119 6885 20131 6919
rect 24946 6916 24952 6928
rect 24907 6888 24952 6916
rect 20073 6879 20131 6885
rect 19337 6851 19395 6857
rect 19337 6848 19349 6851
rect 17727 6820 18460 6848
rect 18524 6820 19349 6848
rect 17727 6817 17739 6820
rect 17681 6811 17739 6817
rect 17405 6783 17463 6789
rect 17405 6749 17417 6783
rect 17451 6749 17463 6783
rect 17405 6743 17463 6749
rect 17497 6783 17555 6789
rect 17497 6749 17509 6783
rect 17543 6780 17555 6783
rect 17770 6780 17776 6792
rect 17543 6752 17776 6780
rect 17543 6749 17555 6752
rect 17497 6743 17555 6749
rect 14182 6672 14188 6724
rect 14240 6712 14246 6724
rect 14338 6715 14396 6721
rect 14338 6712 14350 6715
rect 14240 6684 14350 6712
rect 14240 6672 14246 6684
rect 14338 6681 14350 6684
rect 14384 6681 14396 6715
rect 17420 6712 17448 6743
rect 17770 6740 17776 6752
rect 17828 6780 17834 6792
rect 18524 6789 18552 6820
rect 19337 6817 19349 6820
rect 19383 6848 19395 6851
rect 20088 6848 20116 6879
rect 24946 6876 24952 6888
rect 25004 6876 25010 6928
rect 19383 6820 20208 6848
rect 19383 6817 19395 6820
rect 19337 6811 19395 6817
rect 18233 6783 18291 6789
rect 18233 6780 18245 6783
rect 17828 6752 18245 6780
rect 17828 6740 17834 6752
rect 18233 6749 18245 6752
rect 18279 6749 18291 6783
rect 18233 6743 18291 6749
rect 18325 6783 18383 6789
rect 18325 6749 18337 6783
rect 18371 6749 18383 6783
rect 18325 6743 18383 6749
rect 18509 6783 18567 6789
rect 18509 6749 18521 6783
rect 18555 6749 18567 6783
rect 18690 6780 18696 6792
rect 18651 6752 18696 6780
rect 18509 6743 18567 6749
rect 18340 6712 18368 6743
rect 18690 6740 18696 6752
rect 18748 6740 18754 6792
rect 19242 6780 19248 6792
rect 19203 6752 19248 6780
rect 19242 6740 19248 6752
rect 19300 6740 19306 6792
rect 19429 6783 19487 6789
rect 19429 6749 19441 6783
rect 19475 6780 19487 6783
rect 19518 6780 19524 6792
rect 19475 6752 19524 6780
rect 19475 6749 19487 6752
rect 19429 6743 19487 6749
rect 19518 6740 19524 6752
rect 19576 6740 19582 6792
rect 20180 6780 20208 6820
rect 20438 6808 20444 6860
rect 20496 6848 20502 6860
rect 20901 6851 20959 6857
rect 20901 6848 20913 6851
rect 20496 6820 20913 6848
rect 20496 6808 20502 6820
rect 20901 6817 20913 6820
rect 20947 6817 20959 6851
rect 22094 6848 22100 6860
rect 20901 6811 20959 6817
rect 22066 6808 22100 6848
rect 22152 6848 22158 6860
rect 22189 6851 22247 6857
rect 22189 6848 22201 6851
rect 22152 6820 22201 6848
rect 22152 6808 22158 6820
rect 22189 6817 22201 6820
rect 22235 6817 22247 6851
rect 22189 6811 22247 6817
rect 20806 6780 20812 6792
rect 20180 6752 20812 6780
rect 20806 6740 20812 6752
rect 20864 6740 20870 6792
rect 21082 6780 21088 6792
rect 21043 6752 21088 6780
rect 21082 6740 21088 6752
rect 21140 6740 21146 6792
rect 21266 6780 21272 6792
rect 21227 6752 21272 6780
rect 21266 6740 21272 6752
rect 21324 6740 21330 6792
rect 21361 6783 21419 6789
rect 21361 6749 21373 6783
rect 21407 6780 21419 6783
rect 21821 6783 21879 6789
rect 21407 6752 21772 6780
rect 21407 6749 21419 6752
rect 21361 6743 21419 6749
rect 19702 6712 19708 6724
rect 17420 6684 17540 6712
rect 18340 6684 19708 6712
rect 14338 6675 14396 6681
rect 17512 6656 17540 6684
rect 19702 6672 19708 6684
rect 19760 6672 19766 6724
rect 21634 6712 21640 6724
rect 20180 6684 21128 6712
rect 21595 6684 21640 6712
rect 12434 6644 12440 6656
rect 12084 6616 12440 6644
rect 11885 6607 11943 6613
rect 12434 6604 12440 6616
rect 12492 6604 12498 6656
rect 12802 6644 12808 6656
rect 12763 6616 12808 6644
rect 12802 6604 12808 6616
rect 12860 6604 12866 6656
rect 13541 6647 13599 6653
rect 13541 6613 13553 6647
rect 13587 6644 13599 6647
rect 13998 6644 14004 6656
rect 13587 6616 14004 6644
rect 13587 6613 13599 6616
rect 13541 6607 13599 6613
rect 13998 6604 14004 6616
rect 14056 6604 14062 6656
rect 17126 6644 17132 6656
rect 17087 6616 17132 6644
rect 17126 6604 17132 6616
rect 17184 6604 17190 6656
rect 17494 6644 17500 6656
rect 17407 6616 17500 6644
rect 17494 6604 17500 6616
rect 17552 6644 17558 6656
rect 19978 6644 19984 6656
rect 17552 6616 19984 6644
rect 17552 6604 17558 6616
rect 19978 6604 19984 6616
rect 20036 6604 20042 6656
rect 20180 6653 20208 6684
rect 20165 6647 20223 6653
rect 20165 6613 20177 6647
rect 20211 6613 20223 6647
rect 21100 6644 21128 6684
rect 21634 6672 21640 6684
rect 21692 6672 21698 6724
rect 21744 6712 21772 6752
rect 21821 6749 21833 6783
rect 21867 6780 21879 6783
rect 22066 6780 22094 6808
rect 21867 6752 22094 6780
rect 22649 6783 22707 6789
rect 21867 6749 21879 6752
rect 21821 6743 21879 6749
rect 22649 6749 22661 6783
rect 22695 6780 22707 6783
rect 25225 6783 25283 6789
rect 25225 6780 25237 6783
rect 22695 6752 25237 6780
rect 22695 6749 22707 6752
rect 22649 6743 22707 6749
rect 23584 6724 23612 6752
rect 25225 6749 25237 6752
rect 25271 6749 25283 6783
rect 25225 6743 25283 6749
rect 22002 6712 22008 6724
rect 21744 6684 22008 6712
rect 22002 6672 22008 6684
rect 22060 6672 22066 6724
rect 22922 6721 22928 6724
rect 22916 6712 22928 6721
rect 22883 6684 22928 6712
rect 22916 6675 22928 6684
rect 22922 6672 22928 6675
rect 22980 6672 22986 6724
rect 23566 6672 23572 6724
rect 23624 6672 23630 6724
rect 24670 6672 24676 6724
rect 24728 6712 24734 6724
rect 24765 6715 24823 6721
rect 24765 6712 24777 6715
rect 24728 6684 24777 6712
rect 24728 6672 24734 6684
rect 24765 6681 24777 6684
rect 24811 6681 24823 6715
rect 24765 6675 24823 6681
rect 25492 6715 25550 6721
rect 25492 6681 25504 6715
rect 25538 6712 25550 6715
rect 25682 6712 25688 6724
rect 25538 6684 25688 6712
rect 25538 6681 25550 6684
rect 25492 6675 25550 6681
rect 25682 6672 25688 6684
rect 25740 6672 25746 6724
rect 23382 6644 23388 6656
rect 21100 6616 23388 6644
rect 20165 6607 20223 6613
rect 23382 6604 23388 6616
rect 23440 6604 23446 6656
rect 25130 6604 25136 6656
rect 25188 6644 25194 6656
rect 26605 6647 26663 6653
rect 26605 6644 26617 6647
rect 25188 6616 26617 6644
rect 25188 6604 25194 6616
rect 26605 6613 26617 6616
rect 26651 6613 26663 6647
rect 26605 6607 26663 6613
rect 1104 6554 28888 6576
rect 1104 6502 10214 6554
rect 10266 6502 10278 6554
rect 10330 6502 10342 6554
rect 10394 6502 10406 6554
rect 10458 6502 10470 6554
rect 10522 6502 19478 6554
rect 19530 6502 19542 6554
rect 19594 6502 19606 6554
rect 19658 6502 19670 6554
rect 19722 6502 19734 6554
rect 19786 6502 28888 6554
rect 1104 6480 28888 6502
rect 6362 6400 6368 6452
rect 6420 6440 6426 6452
rect 6457 6443 6515 6449
rect 6457 6440 6469 6443
rect 6420 6412 6469 6440
rect 6420 6400 6426 6412
rect 6457 6409 6469 6412
rect 6503 6409 6515 6443
rect 6457 6403 6515 6409
rect 6638 6400 6644 6452
rect 6696 6440 6702 6452
rect 8110 6440 8116 6452
rect 6696 6412 8116 6440
rect 6696 6400 6702 6412
rect 6748 6381 6776 6412
rect 8110 6400 8116 6412
rect 8168 6400 8174 6452
rect 8386 6440 8392 6452
rect 8347 6412 8392 6440
rect 8386 6400 8392 6412
rect 8444 6400 8450 6452
rect 8478 6400 8484 6452
rect 8536 6440 8542 6452
rect 8757 6443 8815 6449
rect 8757 6440 8769 6443
rect 8536 6412 8769 6440
rect 8536 6400 8542 6412
rect 8757 6409 8769 6412
rect 8803 6409 8815 6443
rect 9858 6440 9864 6452
rect 9819 6412 9864 6440
rect 8757 6403 8815 6409
rect 9858 6400 9864 6412
rect 9916 6400 9922 6452
rect 9950 6400 9956 6452
rect 10008 6400 10014 6452
rect 12710 6400 12716 6452
rect 12768 6440 12774 6452
rect 13541 6443 13599 6449
rect 13541 6440 13553 6443
rect 12768 6412 13553 6440
rect 12768 6400 12774 6412
rect 13541 6409 13553 6412
rect 13587 6409 13599 6443
rect 14182 6440 14188 6452
rect 14240 6449 14246 6452
rect 14149 6412 14188 6440
rect 13541 6403 13599 6409
rect 14182 6400 14188 6412
rect 14240 6403 14249 6449
rect 14277 6443 14335 6449
rect 14277 6409 14289 6443
rect 14323 6440 14335 6443
rect 14829 6443 14887 6449
rect 14829 6440 14841 6443
rect 14323 6412 14841 6440
rect 14323 6409 14335 6412
rect 14277 6403 14335 6409
rect 14829 6409 14841 6412
rect 14875 6409 14887 6443
rect 14829 6403 14887 6409
rect 14240 6400 14246 6403
rect 15930 6400 15936 6452
rect 15988 6440 15994 6452
rect 16301 6443 16359 6449
rect 16301 6440 16313 6443
rect 15988 6412 16313 6440
rect 15988 6400 15994 6412
rect 16301 6409 16313 6412
rect 16347 6409 16359 6443
rect 17954 6440 17960 6452
rect 16301 6403 16359 6409
rect 17696 6412 17960 6440
rect 6733 6375 6791 6381
rect 6733 6341 6745 6375
rect 6779 6341 6791 6375
rect 6733 6335 6791 6341
rect 6963 6375 7021 6381
rect 6963 6341 6975 6375
rect 7009 6372 7021 6375
rect 7742 6372 7748 6384
rect 7009 6344 7748 6372
rect 7009 6341 7021 6344
rect 6963 6335 7021 6341
rect 7742 6332 7748 6344
rect 7800 6332 7806 6384
rect 8021 6375 8079 6381
rect 8021 6341 8033 6375
rect 8067 6341 8079 6375
rect 8021 6335 8079 6341
rect 8237 6375 8295 6381
rect 8237 6341 8249 6375
rect 8283 6372 8295 6375
rect 9766 6372 9772 6384
rect 8283 6344 9772 6372
rect 8283 6341 8295 6344
rect 8237 6335 8295 6341
rect 6641 6307 6699 6313
rect 6641 6273 6653 6307
rect 6687 6273 6699 6307
rect 6641 6267 6699 6273
rect 6656 6168 6684 6267
rect 6822 6264 6828 6316
rect 6880 6304 6886 6316
rect 7098 6304 7104 6316
rect 6880 6276 6973 6304
rect 7059 6276 7104 6304
rect 6880 6264 6886 6276
rect 7098 6264 7104 6276
rect 7156 6304 7162 6316
rect 7377 6307 7435 6313
rect 7377 6304 7389 6307
rect 7156 6276 7389 6304
rect 7156 6264 7162 6276
rect 7377 6273 7389 6276
rect 7423 6273 7435 6307
rect 7558 6304 7564 6316
rect 7519 6276 7564 6304
rect 7377 6267 7435 6273
rect 7558 6264 7564 6276
rect 7616 6264 7622 6316
rect 6840 6236 6868 6264
rect 8036 6236 8064 6335
rect 9766 6332 9772 6344
rect 9824 6332 9830 6384
rect 9968 6372 9996 6400
rect 9968 6344 11008 6372
rect 8849 6307 8907 6313
rect 8849 6304 8861 6307
rect 8312 6276 8861 6304
rect 8312 6248 8340 6276
rect 8849 6273 8861 6276
rect 8895 6273 8907 6307
rect 8849 6267 8907 6273
rect 9677 6307 9735 6313
rect 9677 6273 9689 6307
rect 9723 6273 9735 6307
rect 9677 6267 9735 6273
rect 9953 6307 10011 6313
rect 9953 6273 9965 6307
rect 9999 6304 10011 6307
rect 10594 6304 10600 6316
rect 9999 6276 10600 6304
rect 9999 6273 10011 6276
rect 9953 6267 10011 6273
rect 8294 6236 8300 6248
rect 6840 6208 7512 6236
rect 8036 6208 8300 6236
rect 7377 6171 7435 6177
rect 7377 6168 7389 6171
rect 6656 6140 7389 6168
rect 7377 6137 7389 6140
rect 7423 6137 7435 6171
rect 7484 6168 7512 6208
rect 8294 6196 8300 6208
rect 8352 6196 8358 6248
rect 9692 6236 9720 6267
rect 10594 6264 10600 6276
rect 10652 6264 10658 6316
rect 10980 6313 11008 6344
rect 11054 6332 11060 6384
rect 11112 6372 11118 6384
rect 11609 6375 11667 6381
rect 11609 6372 11621 6375
rect 11112 6344 11621 6372
rect 11112 6332 11118 6344
rect 11609 6341 11621 6344
rect 11655 6341 11667 6375
rect 13906 6372 13912 6384
rect 11609 6335 11667 6341
rect 12176 6344 13912 6372
rect 10965 6307 11023 6313
rect 10965 6273 10977 6307
rect 11011 6273 11023 6307
rect 10965 6267 11023 6273
rect 11149 6307 11207 6313
rect 11149 6273 11161 6307
rect 11195 6273 11207 6307
rect 11149 6267 11207 6273
rect 9858 6236 9864 6248
rect 9692 6208 9864 6236
rect 9858 6196 9864 6208
rect 9916 6236 9922 6248
rect 10134 6236 10140 6248
rect 9916 6208 10140 6236
rect 9916 6196 9922 6208
rect 10134 6196 10140 6208
rect 10192 6196 10198 6248
rect 11164 6236 11192 6267
rect 11882 6236 11888 6248
rect 11164 6208 11888 6236
rect 11882 6196 11888 6208
rect 11940 6196 11946 6248
rect 12176 6245 12204 6344
rect 13906 6332 13912 6344
rect 13964 6332 13970 6384
rect 14642 6332 14648 6384
rect 14700 6372 14706 6384
rect 14700 6344 16160 6372
rect 14700 6332 14706 6344
rect 12250 6264 12256 6316
rect 12308 6304 12314 6316
rect 12417 6307 12475 6313
rect 12417 6304 12429 6307
rect 12308 6276 12429 6304
rect 12308 6264 12314 6276
rect 12417 6273 12429 6276
rect 12463 6273 12475 6307
rect 12417 6267 12475 6273
rect 13998 6264 14004 6316
rect 14056 6304 14062 6316
rect 14093 6307 14151 6313
rect 14093 6304 14105 6307
rect 14056 6276 14105 6304
rect 14056 6264 14062 6276
rect 14093 6273 14105 6276
rect 14139 6273 14151 6307
rect 14093 6267 14151 6273
rect 14366 6264 14372 6316
rect 14424 6304 14430 6316
rect 15028 6313 15056 6344
rect 14829 6307 14887 6313
rect 14424 6276 14469 6304
rect 14424 6264 14430 6276
rect 14829 6273 14841 6307
rect 14875 6273 14887 6307
rect 14829 6267 14887 6273
rect 15013 6307 15071 6313
rect 15013 6273 15025 6307
rect 15059 6273 15071 6307
rect 15013 6267 15071 6273
rect 12161 6239 12219 6245
rect 12161 6236 12173 6239
rect 11992 6208 12173 6236
rect 11992 6180 12020 6208
rect 12161 6205 12173 6208
rect 12207 6205 12219 6239
rect 14844 6236 14872 6267
rect 15470 6264 15476 6316
rect 15528 6304 15534 6316
rect 16132 6313 16160 6344
rect 16025 6307 16083 6313
rect 16025 6304 16037 6307
rect 15528 6276 16037 6304
rect 15528 6264 15534 6276
rect 16025 6273 16037 6276
rect 16071 6273 16083 6307
rect 16025 6267 16083 6273
rect 16117 6307 16175 6313
rect 16117 6273 16129 6307
rect 16163 6304 16175 6307
rect 17494 6304 17500 6316
rect 16163 6276 17500 6304
rect 16163 6273 16175 6276
rect 16117 6267 16175 6273
rect 17494 6264 17500 6276
rect 17552 6264 17558 6316
rect 15488 6236 15516 6264
rect 14844 6208 15516 6236
rect 16301 6239 16359 6245
rect 12161 6199 12219 6205
rect 16301 6205 16313 6239
rect 16347 6236 16359 6239
rect 17126 6236 17132 6248
rect 16347 6208 17132 6236
rect 16347 6205 16359 6208
rect 16301 6199 16359 6205
rect 17126 6196 17132 6208
rect 17184 6196 17190 6248
rect 17696 6236 17724 6412
rect 17954 6400 17960 6412
rect 18012 6440 18018 6452
rect 18690 6440 18696 6452
rect 18012 6412 18696 6440
rect 18012 6400 18018 6412
rect 18690 6400 18696 6412
rect 18748 6400 18754 6452
rect 20993 6443 21051 6449
rect 20993 6440 21005 6443
rect 19812 6412 21005 6440
rect 17865 6375 17923 6381
rect 17865 6341 17877 6375
rect 17911 6372 17923 6375
rect 18046 6372 18052 6384
rect 17911 6344 18052 6372
rect 17911 6341 17923 6344
rect 17865 6335 17923 6341
rect 18046 6332 18052 6344
rect 18104 6332 18110 6384
rect 18598 6372 18604 6384
rect 18156 6344 18604 6372
rect 18156 6313 18184 6344
rect 18598 6332 18604 6344
rect 18656 6372 18662 6384
rect 19812 6381 19840 6412
rect 20993 6409 21005 6412
rect 21039 6409 21051 6443
rect 20993 6403 21051 6409
rect 21266 6400 21272 6452
rect 21324 6440 21330 6452
rect 23293 6443 23351 6449
rect 21324 6412 21956 6440
rect 21324 6400 21330 6412
rect 19797 6375 19855 6381
rect 19797 6372 19809 6375
rect 18656 6344 19104 6372
rect 18656 6332 18662 6344
rect 18141 6307 18199 6313
rect 18141 6273 18153 6307
rect 18187 6273 18199 6307
rect 18141 6267 18199 6273
rect 18325 6307 18383 6313
rect 18325 6273 18337 6307
rect 18371 6304 18383 6307
rect 18966 6304 18972 6316
rect 18371 6276 18972 6304
rect 18371 6273 18383 6276
rect 18325 6267 18383 6273
rect 18966 6264 18972 6276
rect 19024 6264 19030 6316
rect 19076 6313 19104 6344
rect 19168 6344 19809 6372
rect 19168 6313 19196 6344
rect 19797 6341 19809 6344
rect 19843 6341 19855 6375
rect 20254 6372 20260 6384
rect 20215 6344 20260 6372
rect 19797 6335 19855 6341
rect 20254 6332 20260 6344
rect 20312 6332 20318 6384
rect 20548 6344 21864 6372
rect 19061 6307 19119 6313
rect 19061 6273 19073 6307
rect 19107 6273 19119 6307
rect 19061 6267 19119 6273
rect 19153 6307 19211 6313
rect 19153 6273 19165 6307
rect 19199 6273 19211 6307
rect 19153 6267 19211 6273
rect 19337 6307 19395 6313
rect 19337 6273 19349 6307
rect 19383 6273 19395 6307
rect 19337 6267 19395 6273
rect 17328 6208 17724 6236
rect 8478 6168 8484 6180
rect 7484 6140 8484 6168
rect 7377 6131 7435 6137
rect 8478 6128 8484 6140
rect 8536 6128 8542 6180
rect 9674 6168 9680 6180
rect 9635 6140 9680 6168
rect 9674 6128 9680 6140
rect 9732 6128 9738 6180
rect 11793 6171 11851 6177
rect 11793 6137 11805 6171
rect 11839 6168 11851 6171
rect 11974 6168 11980 6180
rect 11839 6140 11980 6168
rect 11839 6137 11851 6140
rect 11793 6131 11851 6137
rect 11974 6128 11980 6140
rect 12032 6128 12038 6180
rect 7558 6060 7564 6112
rect 7616 6100 7622 6112
rect 8205 6103 8263 6109
rect 8205 6100 8217 6103
rect 7616 6072 8217 6100
rect 7616 6060 7622 6072
rect 8205 6069 8217 6072
rect 8251 6069 8263 6103
rect 8205 6063 8263 6069
rect 10965 6103 11023 6109
rect 10965 6069 10977 6103
rect 11011 6100 11023 6103
rect 12066 6100 12072 6112
rect 11011 6072 12072 6100
rect 11011 6069 11023 6072
rect 10965 6063 11023 6069
rect 12066 6060 12072 6072
rect 12124 6060 12130 6112
rect 12342 6060 12348 6112
rect 12400 6100 12406 6112
rect 17328 6100 17356 6208
rect 17770 6196 17776 6248
rect 17828 6236 17834 6248
rect 19352 6236 19380 6267
rect 19978 6264 19984 6316
rect 20036 6304 20042 6316
rect 20548 6313 20576 6344
rect 20441 6307 20499 6313
rect 20441 6304 20453 6307
rect 20036 6276 20453 6304
rect 20036 6264 20042 6276
rect 20441 6273 20453 6276
rect 20487 6273 20499 6307
rect 20441 6267 20499 6273
rect 20533 6307 20591 6313
rect 20533 6273 20545 6307
rect 20579 6273 20591 6307
rect 20533 6267 20591 6273
rect 20901 6307 20959 6313
rect 20901 6273 20913 6307
rect 20947 6304 20959 6307
rect 21082 6304 21088 6316
rect 20947 6276 21088 6304
rect 20947 6273 20959 6276
rect 20901 6267 20959 6273
rect 21082 6264 21088 6276
rect 21140 6264 21146 6316
rect 17828 6208 19380 6236
rect 21269 6239 21327 6245
rect 17828 6196 17834 6208
rect 21269 6205 21281 6239
rect 21315 6236 21327 6239
rect 21358 6236 21364 6248
rect 21315 6208 21364 6236
rect 21315 6205 21327 6208
rect 21269 6199 21327 6205
rect 21358 6196 21364 6208
rect 21416 6196 21422 6248
rect 21836 6245 21864 6344
rect 21821 6239 21879 6245
rect 21821 6205 21833 6239
rect 21867 6205 21879 6239
rect 21928 6236 21956 6412
rect 23293 6409 23305 6443
rect 23339 6440 23351 6443
rect 23934 6440 23940 6452
rect 23339 6412 23940 6440
rect 23339 6409 23351 6412
rect 23293 6403 23351 6409
rect 22922 6372 22928 6384
rect 22883 6344 22928 6372
rect 22922 6332 22928 6344
rect 22980 6332 22986 6384
rect 22002 6264 22008 6316
rect 22060 6304 22066 6316
rect 22189 6307 22247 6313
rect 22189 6304 22201 6307
rect 22060 6276 22201 6304
rect 22060 6264 22066 6276
rect 22189 6273 22201 6276
rect 22235 6273 22247 6307
rect 23106 6304 23112 6316
rect 23067 6276 23112 6304
rect 22189 6267 22247 6273
rect 23106 6264 23112 6276
rect 23164 6264 23170 6316
rect 22097 6239 22155 6245
rect 21928 6208 22048 6236
rect 21821 6199 21879 6205
rect 17402 6128 17408 6180
rect 17460 6168 17466 6180
rect 18877 6171 18935 6177
rect 18877 6168 18889 6171
rect 17460 6140 18889 6168
rect 17460 6128 17466 6140
rect 18877 6137 18889 6140
rect 18923 6137 18935 6171
rect 18877 6131 18935 6137
rect 19426 6128 19432 6180
rect 19484 6168 19490 6180
rect 19981 6171 20039 6177
rect 19981 6168 19993 6171
rect 19484 6140 19993 6168
rect 19484 6128 19490 6140
rect 19981 6137 19993 6140
rect 20027 6168 20039 6171
rect 20070 6168 20076 6180
rect 20027 6140 20076 6168
rect 20027 6137 20039 6140
rect 19981 6131 20039 6137
rect 20070 6128 20076 6140
rect 20128 6168 20134 6180
rect 20990 6168 20996 6180
rect 20128 6140 20996 6168
rect 20128 6128 20134 6140
rect 20990 6128 20996 6140
rect 21048 6128 21054 6180
rect 21177 6171 21235 6177
rect 21177 6137 21189 6171
rect 21223 6168 21235 6171
rect 22020 6168 22048 6208
rect 22097 6205 22109 6239
rect 22143 6205 22155 6239
rect 23014 6236 23020 6248
rect 22975 6208 23020 6236
rect 22097 6199 22155 6205
rect 22112 6168 22140 6199
rect 23014 6196 23020 6208
rect 23072 6196 23078 6248
rect 21223 6140 21956 6168
rect 22020 6140 22140 6168
rect 21223 6137 21235 6140
rect 21177 6131 21235 6137
rect 12400 6072 17356 6100
rect 12400 6060 12406 6072
rect 17862 6060 17868 6112
rect 17920 6100 17926 6112
rect 18233 6103 18291 6109
rect 18233 6100 18245 6103
rect 17920 6072 18245 6100
rect 17920 6060 17926 6072
rect 18233 6069 18245 6072
rect 18279 6069 18291 6103
rect 19058 6100 19064 6112
rect 19019 6072 19064 6100
rect 18233 6063 18291 6069
rect 19058 6060 19064 6072
rect 19116 6060 19122 6112
rect 20254 6060 20260 6112
rect 20312 6100 20318 6112
rect 20349 6103 20407 6109
rect 20349 6100 20361 6103
rect 20312 6072 20361 6100
rect 20312 6060 20318 6072
rect 20349 6069 20361 6072
rect 20395 6069 20407 6103
rect 20349 6063 20407 6069
rect 21085 6103 21143 6109
rect 21085 6069 21097 6103
rect 21131 6100 21143 6103
rect 21818 6100 21824 6112
rect 21131 6072 21824 6100
rect 21131 6069 21143 6072
rect 21085 6063 21143 6069
rect 21818 6060 21824 6072
rect 21876 6060 21882 6112
rect 21928 6100 21956 6140
rect 22186 6100 22192 6112
rect 21928 6072 22192 6100
rect 22186 6060 22192 6072
rect 22244 6100 22250 6112
rect 23308 6100 23336 6403
rect 23934 6400 23940 6412
rect 23992 6400 23998 6452
rect 25682 6440 25688 6452
rect 25643 6412 25688 6440
rect 25682 6400 25688 6412
rect 25740 6400 25746 6452
rect 25314 6372 25320 6384
rect 25275 6344 25320 6372
rect 25314 6332 25320 6344
rect 25372 6332 25378 6384
rect 25406 6332 25412 6384
rect 25464 6372 25470 6384
rect 25464 6344 25509 6372
rect 25464 6332 25470 6344
rect 23382 6264 23388 6316
rect 23440 6304 23446 6316
rect 23842 6304 23848 6316
rect 23440 6276 23533 6304
rect 23803 6276 23848 6304
rect 23440 6264 23446 6276
rect 23842 6264 23848 6276
rect 23900 6264 23906 6316
rect 24670 6304 24676 6316
rect 24631 6276 24676 6304
rect 24670 6264 24676 6276
rect 24728 6264 24734 6316
rect 25130 6304 25136 6316
rect 25091 6276 25136 6304
rect 25130 6264 25136 6276
rect 25188 6264 25194 6316
rect 25501 6307 25559 6313
rect 25501 6273 25513 6307
rect 25547 6273 25559 6307
rect 25501 6267 25559 6273
rect 23400 6236 23428 6264
rect 25516 6236 25544 6267
rect 23400 6208 25544 6236
rect 24854 6168 24860 6180
rect 24815 6140 24860 6168
rect 24854 6128 24860 6140
rect 24912 6128 24918 6180
rect 24026 6100 24032 6112
rect 22244 6072 23336 6100
rect 23987 6072 24032 6100
rect 22244 6060 22250 6072
rect 24026 6060 24032 6072
rect 24084 6060 24090 6112
rect 1104 6010 28888 6032
rect 1104 5958 5582 6010
rect 5634 5958 5646 6010
rect 5698 5958 5710 6010
rect 5762 5958 5774 6010
rect 5826 5958 5838 6010
rect 5890 5958 14846 6010
rect 14898 5958 14910 6010
rect 14962 5958 14974 6010
rect 15026 5958 15038 6010
rect 15090 5958 15102 6010
rect 15154 5958 24110 6010
rect 24162 5958 24174 6010
rect 24226 5958 24238 6010
rect 24290 5958 24302 6010
rect 24354 5958 24366 6010
rect 24418 5958 28888 6010
rect 1104 5936 28888 5958
rect 8478 5896 8484 5908
rect 8439 5868 8484 5896
rect 8478 5856 8484 5868
rect 8536 5856 8542 5908
rect 10686 5896 10692 5908
rect 9140 5868 10692 5896
rect 9140 5828 9168 5868
rect 10686 5856 10692 5868
rect 10744 5856 10750 5908
rect 12161 5899 12219 5905
rect 12161 5865 12173 5899
rect 12207 5896 12219 5899
rect 12250 5896 12256 5908
rect 12207 5868 12256 5896
rect 12207 5865 12219 5868
rect 12161 5859 12219 5865
rect 12250 5856 12256 5868
rect 12308 5856 12314 5908
rect 12894 5856 12900 5908
rect 12952 5896 12958 5908
rect 13265 5899 13323 5905
rect 13265 5896 13277 5899
rect 12952 5868 13277 5896
rect 12952 5856 12958 5868
rect 13265 5865 13277 5868
rect 13311 5865 13323 5899
rect 13265 5859 13323 5865
rect 13354 5856 13360 5908
rect 13412 5896 13418 5908
rect 14369 5899 14427 5905
rect 14369 5896 14381 5899
rect 13412 5868 14381 5896
rect 13412 5856 13418 5868
rect 14369 5865 14381 5868
rect 14415 5865 14427 5899
rect 14369 5859 14427 5865
rect 14553 5899 14611 5905
rect 14553 5865 14565 5899
rect 14599 5865 14611 5899
rect 14553 5859 14611 5865
rect 18325 5899 18383 5905
rect 18325 5865 18337 5899
rect 18371 5896 18383 5899
rect 19058 5896 19064 5908
rect 18371 5868 19064 5896
rect 18371 5865 18383 5868
rect 18325 5859 18383 5865
rect 9048 5800 9168 5828
rect 9217 5831 9275 5837
rect 8110 5720 8116 5772
rect 8168 5760 8174 5772
rect 8570 5760 8576 5772
rect 8168 5732 8576 5760
rect 8168 5720 8174 5732
rect 8570 5720 8576 5732
rect 8628 5720 8634 5772
rect 1673 5695 1731 5701
rect 1673 5661 1685 5695
rect 1719 5692 1731 5695
rect 7857 5695 7915 5701
rect 1719 5664 2774 5692
rect 1719 5661 1731 5664
rect 1673 5655 1731 5661
rect 1486 5556 1492 5568
rect 1447 5528 1492 5556
rect 1486 5516 1492 5528
rect 1544 5516 1550 5568
rect 2746 5556 2774 5664
rect 7857 5661 7869 5695
rect 7903 5692 7915 5695
rect 8478 5692 8484 5704
rect 7903 5664 8484 5692
rect 7903 5661 7915 5664
rect 7857 5655 7915 5661
rect 8478 5652 8484 5664
rect 8536 5652 8542 5704
rect 9048 5701 9076 5800
rect 9217 5797 9229 5831
rect 9263 5828 9275 5831
rect 9674 5828 9680 5840
rect 9263 5800 9680 5828
rect 9263 5797 9275 5800
rect 9217 5791 9275 5797
rect 9674 5788 9680 5800
rect 9732 5788 9738 5840
rect 12342 5828 12348 5840
rect 9784 5800 12348 5828
rect 9306 5760 9312 5772
rect 9267 5732 9312 5760
rect 9306 5720 9312 5732
rect 9364 5720 9370 5772
rect 9784 5701 9812 5800
rect 12342 5788 12348 5800
rect 12400 5788 12406 5840
rect 12526 5788 12532 5840
rect 12584 5828 12590 5840
rect 12710 5828 12716 5840
rect 12584 5800 12716 5828
rect 12584 5788 12590 5800
rect 12710 5788 12716 5800
rect 12768 5828 12774 5840
rect 14568 5828 14596 5859
rect 19058 5856 19064 5868
rect 19116 5856 19122 5908
rect 19426 5896 19432 5908
rect 19387 5868 19432 5896
rect 19426 5856 19432 5868
rect 19484 5856 19490 5908
rect 21266 5856 21272 5908
rect 21324 5896 21330 5908
rect 21729 5899 21787 5905
rect 21729 5896 21741 5899
rect 21324 5868 21741 5896
rect 21324 5856 21330 5868
rect 21729 5865 21741 5868
rect 21775 5865 21787 5899
rect 22186 5896 22192 5908
rect 22147 5868 22192 5896
rect 21729 5859 21787 5865
rect 22186 5856 22192 5868
rect 22244 5856 22250 5908
rect 22465 5899 22523 5905
rect 22465 5865 22477 5899
rect 22511 5865 22523 5899
rect 22465 5859 22523 5865
rect 23569 5899 23627 5905
rect 23569 5865 23581 5899
rect 23615 5896 23627 5899
rect 23842 5896 23848 5908
rect 23615 5868 23848 5896
rect 23615 5865 23627 5868
rect 23569 5859 23627 5865
rect 12768 5800 14596 5828
rect 14921 5831 14979 5837
rect 12768 5788 12774 5800
rect 14921 5797 14933 5831
rect 14967 5828 14979 5831
rect 15378 5828 15384 5840
rect 14967 5800 15384 5828
rect 14967 5797 14979 5800
rect 14921 5791 14979 5797
rect 15378 5788 15384 5800
rect 15436 5788 15442 5840
rect 16853 5831 16911 5837
rect 16853 5797 16865 5831
rect 16899 5828 16911 5831
rect 16942 5828 16948 5840
rect 16899 5800 16948 5828
rect 16899 5797 16911 5800
rect 16853 5791 16911 5797
rect 16942 5788 16948 5800
rect 17000 5788 17006 5840
rect 18782 5828 18788 5840
rect 17328 5800 18788 5828
rect 10778 5760 10784 5772
rect 9876 5732 10784 5760
rect 9876 5701 9904 5732
rect 10778 5720 10784 5732
rect 10836 5760 10842 5772
rect 10836 5732 11008 5760
rect 10836 5720 10842 5732
rect 9033 5695 9091 5701
rect 9033 5661 9045 5695
rect 9079 5661 9091 5695
rect 9033 5655 9091 5661
rect 9125 5695 9183 5701
rect 9125 5661 9137 5695
rect 9171 5692 9183 5695
rect 9769 5695 9827 5701
rect 9171 5664 9720 5692
rect 9171 5661 9183 5664
rect 9125 5655 9183 5661
rect 6733 5559 6791 5565
rect 6733 5556 6745 5559
rect 2746 5528 6745 5556
rect 6733 5525 6745 5528
rect 6779 5525 6791 5559
rect 9582 5556 9588 5568
rect 9543 5528 9588 5556
rect 6733 5519 6791 5525
rect 9582 5516 9588 5528
rect 9640 5516 9646 5568
rect 9692 5556 9720 5664
rect 9769 5661 9781 5695
rect 9815 5661 9827 5695
rect 9769 5655 9827 5661
rect 9861 5695 9919 5701
rect 9861 5661 9873 5695
rect 9907 5661 9919 5695
rect 10042 5692 10048 5704
rect 10003 5664 10048 5692
rect 9861 5655 9919 5661
rect 10042 5652 10048 5664
rect 10100 5652 10106 5704
rect 10134 5652 10140 5704
rect 10192 5692 10198 5704
rect 10192 5664 10237 5692
rect 10192 5652 10198 5664
rect 10594 5652 10600 5704
rect 10652 5692 10658 5704
rect 10980 5701 11008 5732
rect 13170 5720 13176 5772
rect 13228 5760 13234 5772
rect 13357 5763 13415 5769
rect 13357 5760 13369 5763
rect 13228 5732 13369 5760
rect 13228 5720 13234 5732
rect 13357 5729 13369 5732
rect 13403 5729 13415 5763
rect 13357 5723 13415 5729
rect 10865 5695 10923 5701
rect 10865 5692 10877 5695
rect 10652 5664 10877 5692
rect 10652 5652 10658 5664
rect 10865 5661 10877 5664
rect 10911 5661 10923 5695
rect 10865 5655 10923 5661
rect 10957 5695 11015 5701
rect 10957 5661 10969 5695
rect 11003 5661 11015 5695
rect 11149 5695 11207 5701
rect 11149 5692 11161 5695
rect 10957 5655 11015 5661
rect 11072 5664 11161 5692
rect 11072 5636 11100 5664
rect 11149 5661 11161 5664
rect 11195 5661 11207 5695
rect 11149 5655 11207 5661
rect 11251 5695 11309 5701
rect 11251 5661 11263 5695
rect 11297 5692 11309 5695
rect 11514 5692 11520 5704
rect 11297 5664 11376 5692
rect 11475 5664 11520 5692
rect 11297 5661 11309 5664
rect 11251 5655 11309 5661
rect 11054 5584 11060 5636
rect 11112 5584 11118 5636
rect 11348 5624 11376 5664
rect 11514 5652 11520 5664
rect 11572 5652 11578 5704
rect 11698 5692 11704 5704
rect 11659 5664 11704 5692
rect 11698 5652 11704 5664
rect 11756 5652 11762 5704
rect 11790 5652 11796 5704
rect 11848 5692 11854 5704
rect 11931 5695 11989 5701
rect 11848 5664 11893 5692
rect 11848 5652 11854 5664
rect 11931 5661 11943 5695
rect 11977 5692 11989 5695
rect 12066 5692 12072 5704
rect 11977 5664 12072 5692
rect 11977 5661 11989 5664
rect 11931 5655 11989 5661
rect 12066 5652 12072 5664
rect 12124 5652 12130 5704
rect 12434 5652 12440 5704
rect 12492 5692 12498 5704
rect 13541 5695 13599 5701
rect 13541 5692 13553 5695
rect 12492 5664 13553 5692
rect 12492 5652 12498 5664
rect 13541 5661 13553 5664
rect 13587 5692 13599 5695
rect 13906 5692 13912 5704
rect 13587 5664 13912 5692
rect 13587 5661 13599 5664
rect 13541 5655 13599 5661
rect 13906 5652 13912 5664
rect 13964 5652 13970 5704
rect 16574 5692 16580 5704
rect 16535 5664 16580 5692
rect 16574 5652 16580 5664
rect 16632 5652 16638 5704
rect 16669 5695 16727 5701
rect 16669 5661 16681 5695
rect 16715 5692 16727 5695
rect 17328 5692 17356 5800
rect 18782 5788 18788 5800
rect 18840 5788 18846 5840
rect 17770 5720 17776 5772
rect 17828 5760 17834 5772
rect 18141 5763 18199 5769
rect 18141 5760 18153 5763
rect 17828 5732 18153 5760
rect 17828 5720 17834 5732
rect 18141 5729 18153 5732
rect 18187 5760 18199 5763
rect 19076 5760 19104 5856
rect 21361 5831 21419 5837
rect 21361 5797 21373 5831
rect 21407 5828 21419 5831
rect 21818 5828 21824 5840
rect 21407 5800 21824 5828
rect 21407 5797 21419 5800
rect 21361 5791 21419 5797
rect 21818 5788 21824 5800
rect 21876 5788 21882 5840
rect 19337 5763 19395 5769
rect 19337 5760 19349 5763
rect 18187 5732 18460 5760
rect 19076 5732 19349 5760
rect 18187 5729 18199 5732
rect 18141 5723 18199 5729
rect 16715 5664 17356 5692
rect 17405 5695 17463 5701
rect 16715 5661 16727 5664
rect 16669 5655 16727 5661
rect 17405 5661 17417 5695
rect 17451 5661 17463 5695
rect 17405 5655 17463 5661
rect 17681 5695 17739 5701
rect 17681 5661 17693 5695
rect 17727 5692 17739 5695
rect 17862 5692 17868 5704
rect 17727 5664 17868 5692
rect 17727 5661 17739 5664
rect 17681 5655 17739 5661
rect 12158 5624 12164 5636
rect 11348 5596 12164 5624
rect 12158 5584 12164 5596
rect 12216 5584 12222 5636
rect 12621 5627 12679 5633
rect 12621 5593 12633 5627
rect 12667 5593 12679 5627
rect 13078 5624 13084 5636
rect 12621 5587 12679 5593
rect 12820 5596 13084 5624
rect 9950 5556 9956 5568
rect 9692 5528 9956 5556
rect 9950 5516 9956 5528
rect 10008 5516 10014 5568
rect 10686 5556 10692 5568
rect 10647 5528 10692 5556
rect 10686 5516 10692 5528
rect 10744 5516 10750 5568
rect 11330 5516 11336 5568
rect 11388 5556 11394 5568
rect 11790 5556 11796 5568
rect 11388 5528 11796 5556
rect 11388 5516 11394 5528
rect 11790 5516 11796 5528
rect 11848 5556 11854 5568
rect 12529 5559 12587 5565
rect 12529 5556 12541 5559
rect 11848 5528 12541 5556
rect 11848 5516 11854 5528
rect 12529 5525 12541 5528
rect 12575 5525 12587 5559
rect 12636 5556 12664 5587
rect 12820 5556 12848 5596
rect 13078 5584 13084 5596
rect 13136 5584 13142 5636
rect 13265 5627 13323 5633
rect 13265 5593 13277 5627
rect 13311 5624 13323 5627
rect 13354 5624 13360 5636
rect 13311 5596 13360 5624
rect 13311 5593 13323 5596
rect 13265 5587 13323 5593
rect 13354 5584 13360 5596
rect 13412 5584 13418 5636
rect 14550 5624 14556 5636
rect 14511 5596 14556 5624
rect 14550 5584 14556 5596
rect 14608 5584 14614 5636
rect 16853 5627 16911 5633
rect 16853 5593 16865 5627
rect 16899 5624 16911 5627
rect 17221 5627 17279 5633
rect 17221 5624 17233 5627
rect 16899 5596 17233 5624
rect 16899 5593 16911 5596
rect 16853 5587 16911 5593
rect 17221 5593 17233 5596
rect 17267 5593 17279 5627
rect 17420 5624 17448 5655
rect 17862 5652 17868 5664
rect 17920 5652 17926 5704
rect 17954 5652 17960 5704
rect 18012 5652 18018 5704
rect 18322 5692 18328 5704
rect 18283 5664 18328 5692
rect 18322 5652 18328 5664
rect 18380 5652 18386 5704
rect 18432 5692 18460 5732
rect 19337 5729 19349 5732
rect 19383 5729 19395 5763
rect 19337 5723 19395 5729
rect 19886 5720 19892 5772
rect 19944 5760 19950 5772
rect 19981 5763 20039 5769
rect 19981 5760 19993 5763
rect 19944 5732 19993 5760
rect 19944 5720 19950 5732
rect 19981 5729 19993 5732
rect 20027 5729 20039 5763
rect 19981 5723 20039 5729
rect 20990 5720 20996 5772
rect 21048 5760 21054 5772
rect 22480 5760 22508 5859
rect 23842 5856 23848 5868
rect 23900 5856 23906 5908
rect 22833 5831 22891 5837
rect 22833 5797 22845 5831
rect 22879 5797 22891 5831
rect 22833 5791 22891 5797
rect 23293 5831 23351 5837
rect 23293 5797 23305 5831
rect 23339 5828 23351 5831
rect 23750 5828 23756 5840
rect 23339 5800 23756 5828
rect 23339 5797 23351 5800
rect 23293 5791 23351 5797
rect 21048 5732 22508 5760
rect 22848 5760 22876 5791
rect 23750 5788 23756 5800
rect 23808 5788 23814 5840
rect 24670 5760 24676 5772
rect 22848 5732 24676 5760
rect 21048 5720 21054 5732
rect 24670 5720 24676 5732
rect 24728 5760 24734 5772
rect 24949 5763 25007 5769
rect 24949 5760 24961 5763
rect 24728 5732 24961 5760
rect 24728 5720 24734 5732
rect 24949 5729 24961 5732
rect 24995 5729 25007 5763
rect 24949 5723 25007 5729
rect 20254 5701 20260 5704
rect 19245 5695 19303 5701
rect 19245 5692 19257 5695
rect 18432 5664 19257 5692
rect 19245 5661 19257 5664
rect 19291 5661 19303 5695
rect 20248 5692 20260 5701
rect 20215 5664 20260 5692
rect 19245 5655 19303 5661
rect 20248 5655 20260 5664
rect 20254 5652 20260 5655
rect 20312 5652 20318 5704
rect 21358 5652 21364 5704
rect 21416 5692 21422 5704
rect 21913 5695 21971 5701
rect 21913 5692 21925 5695
rect 21416 5664 21925 5692
rect 21416 5652 21422 5664
rect 21913 5661 21925 5664
rect 21959 5661 21971 5695
rect 21913 5655 21971 5661
rect 22005 5695 22063 5701
rect 22005 5661 22017 5695
rect 22051 5692 22063 5695
rect 22094 5692 22100 5704
rect 22051 5664 22100 5692
rect 22051 5661 22063 5664
rect 22005 5655 22063 5661
rect 22094 5652 22100 5664
rect 22152 5652 22158 5704
rect 22465 5695 22523 5701
rect 22465 5692 22477 5695
rect 22204 5664 22477 5692
rect 17972 5624 18000 5652
rect 17420 5596 18000 5624
rect 18049 5627 18107 5633
rect 17221 5587 17279 5593
rect 18049 5593 18061 5627
rect 18095 5624 18107 5627
rect 18138 5624 18144 5636
rect 18095 5596 18144 5624
rect 18095 5593 18107 5596
rect 18049 5587 18107 5593
rect 18138 5584 18144 5596
rect 18196 5584 18202 5636
rect 19334 5624 19340 5636
rect 18524 5596 19340 5624
rect 12636 5528 12848 5556
rect 13725 5559 13783 5565
rect 12529 5519 12587 5525
rect 13725 5525 13737 5559
rect 13771 5556 13783 5559
rect 14274 5556 14280 5568
rect 13771 5528 14280 5556
rect 13771 5525 13783 5528
rect 13725 5519 13783 5525
rect 14274 5516 14280 5528
rect 14332 5516 14338 5568
rect 17402 5516 17408 5568
rect 17460 5556 17466 5568
rect 17589 5559 17647 5565
rect 17589 5556 17601 5559
rect 17460 5528 17601 5556
rect 17460 5516 17466 5528
rect 17589 5525 17601 5528
rect 17635 5525 17647 5559
rect 17589 5519 17647 5525
rect 17862 5516 17868 5568
rect 17920 5556 17926 5568
rect 18524 5565 18552 5596
rect 19334 5584 19340 5596
rect 19392 5624 19398 5636
rect 22204 5633 22232 5664
rect 22465 5661 22477 5664
rect 22511 5661 22523 5695
rect 22646 5692 22652 5704
rect 22607 5664 22652 5692
rect 22465 5655 22523 5661
rect 22646 5652 22652 5664
rect 22704 5652 22710 5704
rect 23750 5692 23756 5704
rect 23711 5664 23756 5692
rect 23750 5652 23756 5664
rect 23808 5652 23814 5704
rect 24765 5695 24823 5701
rect 24765 5661 24777 5695
rect 24811 5692 24823 5695
rect 25130 5692 25136 5704
rect 24811 5664 25136 5692
rect 24811 5661 24823 5664
rect 24765 5655 24823 5661
rect 25130 5652 25136 5664
rect 25188 5652 25194 5704
rect 28350 5692 28356 5704
rect 28311 5664 28356 5692
rect 28350 5652 28356 5664
rect 28408 5652 28414 5704
rect 22189 5627 22247 5633
rect 22189 5624 22201 5627
rect 19392 5596 22201 5624
rect 19392 5584 19398 5596
rect 22189 5593 22201 5596
rect 22235 5593 22247 5627
rect 22189 5587 22247 5593
rect 23937 5627 23995 5633
rect 23937 5593 23949 5627
rect 23983 5593 23995 5627
rect 23937 5587 23995 5593
rect 18509 5559 18567 5565
rect 18509 5556 18521 5559
rect 17920 5528 18521 5556
rect 17920 5516 17926 5528
rect 18509 5525 18521 5528
rect 18555 5525 18567 5559
rect 18509 5519 18567 5525
rect 18966 5516 18972 5568
rect 19024 5556 19030 5568
rect 19613 5559 19671 5565
rect 19613 5556 19625 5559
rect 19024 5528 19625 5556
rect 19024 5516 19030 5528
rect 19613 5525 19625 5528
rect 19659 5525 19671 5559
rect 19613 5519 19671 5525
rect 20346 5516 20352 5568
rect 20404 5556 20410 5568
rect 22554 5556 22560 5568
rect 20404 5528 22560 5556
rect 20404 5516 20410 5528
rect 22554 5516 22560 5528
rect 22612 5556 22618 5568
rect 23014 5556 23020 5568
rect 22612 5528 23020 5556
rect 22612 5516 22618 5528
rect 23014 5516 23020 5528
rect 23072 5516 23078 5568
rect 23952 5556 23980 5587
rect 24397 5559 24455 5565
rect 24397 5556 24409 5559
rect 23952 5528 24409 5556
rect 24397 5525 24409 5528
rect 24443 5525 24455 5559
rect 24397 5519 24455 5525
rect 24857 5559 24915 5565
rect 24857 5525 24869 5559
rect 24903 5556 24915 5559
rect 25222 5556 25228 5568
rect 24903 5528 25228 5556
rect 24903 5525 24915 5528
rect 24857 5519 24915 5525
rect 25222 5516 25228 5528
rect 25280 5516 25286 5568
rect 1104 5466 28888 5488
rect 1104 5414 10214 5466
rect 10266 5414 10278 5466
rect 10330 5414 10342 5466
rect 10394 5414 10406 5466
rect 10458 5414 10470 5466
rect 10522 5414 19478 5466
rect 19530 5414 19542 5466
rect 19594 5414 19606 5466
rect 19658 5414 19670 5466
rect 19722 5414 19734 5466
rect 19786 5414 28888 5466
rect 1104 5392 28888 5414
rect 9306 5352 9312 5364
rect 9267 5324 9312 5352
rect 9306 5312 9312 5324
rect 9364 5312 9370 5364
rect 9674 5352 9680 5364
rect 9635 5324 9680 5352
rect 9674 5312 9680 5324
rect 9732 5312 9738 5364
rect 11238 5352 11244 5364
rect 10244 5324 11244 5352
rect 8110 5244 8116 5296
rect 8168 5244 8174 5296
rect 9858 5284 9864 5296
rect 9819 5256 9864 5284
rect 9858 5244 9864 5256
rect 9916 5244 9922 5296
rect 7929 5219 7987 5225
rect 7929 5185 7941 5219
rect 7975 5216 7987 5219
rect 8128 5216 8156 5244
rect 7975 5188 8156 5216
rect 8196 5219 8254 5225
rect 7975 5185 7987 5188
rect 7929 5179 7987 5185
rect 8196 5185 8208 5219
rect 8242 5216 8254 5219
rect 9582 5216 9588 5228
rect 8242 5188 9076 5216
rect 9543 5188 9588 5216
rect 8242 5185 8254 5188
rect 8196 5179 8254 5185
rect 9048 5080 9076 5188
rect 9582 5176 9588 5188
rect 9640 5176 9646 5228
rect 10134 5216 10140 5228
rect 10095 5188 10140 5216
rect 10134 5176 10140 5188
rect 10192 5176 10198 5228
rect 10244 5225 10272 5324
rect 11238 5312 11244 5324
rect 11296 5312 11302 5364
rect 11514 5352 11520 5364
rect 11475 5324 11520 5352
rect 11514 5312 11520 5324
rect 11572 5312 11578 5364
rect 11882 5312 11888 5364
rect 11940 5352 11946 5364
rect 12345 5355 12403 5361
rect 12345 5352 12357 5355
rect 11940 5324 12357 5352
rect 11940 5312 11946 5324
rect 12345 5321 12357 5324
rect 12391 5321 12403 5355
rect 12345 5315 12403 5321
rect 16114 5312 16120 5364
rect 16172 5312 16178 5364
rect 17862 5352 17868 5364
rect 16592 5324 17868 5352
rect 10413 5287 10471 5293
rect 10413 5253 10425 5287
rect 10459 5284 10471 5287
rect 10781 5287 10839 5293
rect 10781 5284 10793 5287
rect 10459 5256 10793 5284
rect 10459 5253 10471 5256
rect 10413 5247 10471 5253
rect 10781 5253 10793 5256
rect 10827 5253 10839 5287
rect 11256 5284 11284 5312
rect 12250 5284 12256 5296
rect 11256 5256 12256 5284
rect 10781 5247 10839 5253
rect 12250 5244 12256 5256
rect 12308 5244 12314 5296
rect 13909 5287 13967 5293
rect 12912 5256 13676 5284
rect 12912 5228 12940 5256
rect 10229 5219 10287 5225
rect 10229 5185 10241 5219
rect 10275 5185 10287 5219
rect 10686 5216 10692 5228
rect 10647 5188 10692 5216
rect 10229 5179 10287 5185
rect 10686 5176 10692 5188
rect 10744 5176 10750 5228
rect 10870 5176 10876 5228
rect 10928 5216 10934 5228
rect 10965 5219 11023 5225
rect 10965 5216 10977 5219
rect 10928 5188 10977 5216
rect 10928 5176 10934 5188
rect 10965 5185 10977 5188
rect 11011 5185 11023 5219
rect 11790 5216 11796 5228
rect 11751 5188 11796 5216
rect 10965 5179 11023 5185
rect 11790 5176 11796 5188
rect 11848 5176 11854 5228
rect 12069 5219 12127 5225
rect 12069 5185 12081 5219
rect 12115 5185 12127 5219
rect 12069 5179 12127 5185
rect 10410 5148 10416 5160
rect 10371 5120 10416 5148
rect 10410 5108 10416 5120
rect 10468 5108 10474 5160
rect 9861 5083 9919 5089
rect 9861 5080 9873 5083
rect 9048 5052 9873 5080
rect 9861 5049 9873 5052
rect 9907 5049 9919 5083
rect 9861 5043 9919 5049
rect 9950 5040 9956 5092
rect 10008 5080 10014 5092
rect 10965 5083 11023 5089
rect 10965 5080 10977 5083
rect 10008 5052 10977 5080
rect 10008 5040 10014 5052
rect 10965 5049 10977 5052
rect 11011 5049 11023 5083
rect 12084 5080 12112 5179
rect 12158 5176 12164 5228
rect 12216 5216 12222 5228
rect 12713 5219 12771 5225
rect 12713 5216 12725 5219
rect 12216 5188 12725 5216
rect 12216 5176 12222 5188
rect 12713 5185 12725 5188
rect 12759 5216 12771 5219
rect 12894 5216 12900 5228
rect 12759 5188 12900 5216
rect 12759 5185 12771 5188
rect 12713 5179 12771 5185
rect 12894 5176 12900 5188
rect 12952 5176 12958 5228
rect 12989 5219 13047 5225
rect 12989 5185 13001 5219
rect 13035 5216 13047 5219
rect 13354 5216 13360 5228
rect 13035 5188 13360 5216
rect 13035 5185 13047 5188
rect 12989 5179 13047 5185
rect 13354 5176 13360 5188
rect 13412 5176 13418 5228
rect 13648 5225 13676 5256
rect 13909 5253 13921 5287
rect 13955 5284 13967 5287
rect 14369 5287 14427 5293
rect 14369 5284 14381 5287
rect 13955 5256 14381 5284
rect 13955 5253 13967 5256
rect 13909 5247 13967 5253
rect 14369 5253 14381 5256
rect 14415 5253 14427 5287
rect 15286 5284 15292 5296
rect 14369 5247 14427 5253
rect 15120 5256 15292 5284
rect 13633 5219 13691 5225
rect 13633 5185 13645 5219
rect 13679 5185 13691 5219
rect 13633 5179 13691 5185
rect 13998 5176 14004 5228
rect 14056 5216 14062 5228
rect 14185 5219 14243 5225
rect 14185 5216 14197 5219
rect 14056 5188 14197 5216
rect 14056 5176 14062 5188
rect 14185 5185 14197 5188
rect 14231 5185 14243 5219
rect 14185 5179 14243 5185
rect 14274 5176 14280 5228
rect 14332 5216 14338 5228
rect 15120 5225 15148 5256
rect 15286 5244 15292 5256
rect 15344 5284 15350 5296
rect 16132 5284 16160 5312
rect 15344 5256 16160 5284
rect 15344 5244 15350 5256
rect 14461 5219 14519 5225
rect 14461 5216 14473 5219
rect 14332 5188 14473 5216
rect 14332 5176 14338 5188
rect 14461 5185 14473 5188
rect 14507 5185 14519 5219
rect 14461 5179 14519 5185
rect 15105 5219 15163 5225
rect 15105 5185 15117 5219
rect 15151 5185 15163 5219
rect 15105 5179 15163 5185
rect 15657 5219 15715 5225
rect 15657 5185 15669 5219
rect 15703 5185 15715 5219
rect 16117 5219 16175 5225
rect 16117 5216 16129 5219
rect 15657 5179 15715 5185
rect 15948 5188 16129 5216
rect 12618 5148 12624 5160
rect 12579 5120 12624 5148
rect 12618 5108 12624 5120
rect 12676 5108 12682 5160
rect 13078 5148 13084 5160
rect 13039 5120 13084 5148
rect 13078 5108 13084 5120
rect 13136 5108 13142 5160
rect 13906 5148 13912 5160
rect 13867 5120 13912 5148
rect 13906 5108 13912 5120
rect 13964 5108 13970 5160
rect 14550 5108 14556 5160
rect 14608 5148 14614 5160
rect 15013 5151 15071 5157
rect 15013 5148 15025 5151
rect 14608 5120 15025 5148
rect 14608 5108 14614 5120
rect 15013 5117 15025 5120
rect 15059 5148 15071 5151
rect 15672 5148 15700 5179
rect 15059 5120 15700 5148
rect 15059 5117 15071 5120
rect 15013 5111 15071 5117
rect 15948 5080 15976 5188
rect 16117 5185 16129 5188
rect 16163 5185 16175 5219
rect 16117 5179 16175 5185
rect 16025 5151 16083 5157
rect 16025 5117 16037 5151
rect 16071 5148 16083 5151
rect 16592 5148 16620 5324
rect 17862 5312 17868 5324
rect 17920 5312 17926 5364
rect 18049 5355 18107 5361
rect 18049 5321 18061 5355
rect 18095 5352 18107 5355
rect 18322 5352 18328 5364
rect 18095 5324 18328 5352
rect 18095 5321 18107 5324
rect 18049 5315 18107 5321
rect 18322 5312 18328 5324
rect 18380 5312 18386 5364
rect 19613 5355 19671 5361
rect 19613 5321 19625 5355
rect 19659 5352 19671 5355
rect 19886 5352 19892 5364
rect 19659 5324 19892 5352
rect 19659 5321 19671 5324
rect 19613 5315 19671 5321
rect 19886 5312 19892 5324
rect 19944 5312 19950 5364
rect 22002 5352 22008 5364
rect 21744 5324 22008 5352
rect 16758 5284 16764 5296
rect 16671 5256 16764 5284
rect 16684 5225 16712 5256
rect 16758 5244 16764 5256
rect 16816 5284 16822 5296
rect 17586 5284 17592 5296
rect 16816 5256 17592 5284
rect 16816 5244 16822 5256
rect 17586 5244 17592 5256
rect 17644 5244 17650 5296
rect 19705 5287 19763 5293
rect 19705 5253 19717 5287
rect 19751 5284 19763 5287
rect 21634 5284 21640 5296
rect 19751 5256 21640 5284
rect 19751 5253 19763 5256
rect 19705 5247 19763 5253
rect 21634 5244 21640 5256
rect 21692 5244 21698 5296
rect 16942 5225 16948 5228
rect 16669 5219 16727 5225
rect 16669 5185 16681 5219
rect 16715 5185 16727 5219
rect 16936 5216 16948 5225
rect 16903 5188 16948 5216
rect 16669 5179 16727 5185
rect 16936 5179 16948 5188
rect 16942 5176 16948 5179
rect 17000 5176 17006 5228
rect 18322 5216 18328 5228
rect 18283 5188 18328 5216
rect 18322 5176 18328 5188
rect 18380 5176 18386 5228
rect 18598 5216 18604 5228
rect 18559 5188 18604 5216
rect 18598 5176 18604 5188
rect 18656 5176 18662 5228
rect 19242 5176 19248 5228
rect 19300 5216 19306 5228
rect 21744 5216 21772 5324
rect 22002 5312 22008 5324
rect 22060 5352 22066 5364
rect 22741 5355 22799 5361
rect 22741 5352 22753 5355
rect 22060 5324 22753 5352
rect 22060 5312 22066 5324
rect 22741 5321 22753 5324
rect 22787 5321 22799 5355
rect 22741 5315 22799 5321
rect 22281 5287 22339 5293
rect 22281 5253 22293 5287
rect 22327 5284 22339 5287
rect 22646 5284 22652 5296
rect 22327 5256 22652 5284
rect 22327 5253 22339 5256
rect 22281 5247 22339 5253
rect 22646 5244 22652 5256
rect 22704 5244 22710 5296
rect 24026 5293 24032 5296
rect 24020 5284 24032 5293
rect 23987 5256 24032 5284
rect 24020 5247 24032 5256
rect 24026 5244 24032 5247
rect 24084 5244 24090 5296
rect 21910 5216 21916 5228
rect 19300 5188 21772 5216
rect 21871 5188 21916 5216
rect 19300 5176 19306 5188
rect 21910 5176 21916 5188
rect 21968 5176 21974 5228
rect 22097 5219 22155 5225
rect 22097 5185 22109 5219
rect 22143 5185 22155 5219
rect 22097 5179 22155 5185
rect 16071 5120 16620 5148
rect 16071 5117 16083 5120
rect 16025 5111 16083 5117
rect 21542 5108 21548 5160
rect 21600 5148 21606 5160
rect 22112 5148 22140 5179
rect 23014 5176 23020 5228
rect 23072 5216 23078 5228
rect 23109 5219 23167 5225
rect 23109 5216 23121 5219
rect 23072 5188 23121 5216
rect 23072 5176 23078 5188
rect 23109 5185 23121 5188
rect 23155 5185 23167 5219
rect 23109 5179 23167 5185
rect 23293 5219 23351 5225
rect 23293 5185 23305 5219
rect 23339 5216 23351 5219
rect 24854 5216 24860 5228
rect 23339 5188 24860 5216
rect 23339 5185 23351 5188
rect 23293 5179 23351 5185
rect 24854 5176 24860 5188
rect 24912 5176 24918 5228
rect 21600 5120 22140 5148
rect 21600 5108 21606 5120
rect 23566 5108 23572 5160
rect 23624 5148 23630 5160
rect 23753 5151 23811 5157
rect 23753 5148 23765 5151
rect 23624 5120 23765 5148
rect 23624 5108 23630 5120
rect 23753 5117 23765 5120
rect 23799 5117 23811 5151
rect 23753 5111 23811 5117
rect 12084 5052 14780 5080
rect 15948 5052 16712 5080
rect 10965 5043 11023 5049
rect 14752 5024 14780 5052
rect 10042 4972 10048 5024
rect 10100 5012 10106 5024
rect 11054 5012 11060 5024
rect 10100 4984 11060 5012
rect 10100 4972 10106 4984
rect 11054 4972 11060 4984
rect 11112 5012 11118 5024
rect 11698 5012 11704 5024
rect 11112 4984 11704 5012
rect 11112 4972 11118 4984
rect 11698 4972 11704 4984
rect 11756 4972 11762 5024
rect 12434 4972 12440 5024
rect 12492 5012 12498 5024
rect 12529 5015 12587 5021
rect 12529 5012 12541 5015
rect 12492 4984 12541 5012
rect 12492 4972 12498 4984
rect 12529 4981 12541 4984
rect 12575 5012 12587 5015
rect 12894 5012 12900 5024
rect 12575 4984 12900 5012
rect 12575 4981 12587 4984
rect 12529 4975 12587 4981
rect 12894 4972 12900 4984
rect 12952 4972 12958 5024
rect 13170 5012 13176 5024
rect 13131 4984 13176 5012
rect 13170 4972 13176 4984
rect 13228 4972 13234 5024
rect 13357 5015 13415 5021
rect 13357 4981 13369 5015
rect 13403 5012 13415 5015
rect 13446 5012 13452 5024
rect 13403 4984 13452 5012
rect 13403 4981 13415 4984
rect 13357 4975 13415 4981
rect 13446 4972 13452 4984
rect 13504 4972 13510 5024
rect 13538 4972 13544 5024
rect 13596 5012 13602 5024
rect 13725 5015 13783 5021
rect 13725 5012 13737 5015
rect 13596 4984 13737 5012
rect 13596 4972 13602 4984
rect 13725 4981 13737 4984
rect 13771 4981 13783 5015
rect 14182 5012 14188 5024
rect 14143 4984 14188 5012
rect 13725 4975 13783 4981
rect 14182 4972 14188 4984
rect 14240 4972 14246 5024
rect 14734 5012 14740 5024
rect 14695 4984 14740 5012
rect 14734 4972 14740 4984
rect 14792 4972 14798 5024
rect 15378 4972 15384 5024
rect 15436 5012 15442 5024
rect 15749 5015 15807 5021
rect 15749 5012 15761 5015
rect 15436 4984 15761 5012
rect 15436 4972 15442 4984
rect 15749 4981 15761 4984
rect 15795 4981 15807 5015
rect 15749 4975 15807 4981
rect 16114 4972 16120 5024
rect 16172 5012 16178 5024
rect 16301 5015 16359 5021
rect 16301 5012 16313 5015
rect 16172 4984 16313 5012
rect 16172 4972 16178 4984
rect 16301 4981 16313 4984
rect 16347 4981 16359 5015
rect 16684 5012 16712 5052
rect 17954 5012 17960 5024
rect 16684 4984 17960 5012
rect 16301 4975 16359 4981
rect 17954 4972 17960 4984
rect 18012 5012 18018 5024
rect 19242 5012 19248 5024
rect 18012 4984 19248 5012
rect 18012 4972 18018 4984
rect 19242 4972 19248 4984
rect 19300 4972 19306 5024
rect 23106 5012 23112 5024
rect 23067 4984 23112 5012
rect 23106 4972 23112 4984
rect 23164 4972 23170 5024
rect 23768 5012 23796 5111
rect 24486 5012 24492 5024
rect 23768 4984 24492 5012
rect 24486 4972 24492 4984
rect 24544 4972 24550 5024
rect 25133 5015 25191 5021
rect 25133 4981 25145 5015
rect 25179 5012 25191 5015
rect 25222 5012 25228 5024
rect 25179 4984 25228 5012
rect 25179 4981 25191 4984
rect 25133 4975 25191 4981
rect 25222 4972 25228 4984
rect 25280 4972 25286 5024
rect 1104 4922 28888 4944
rect 1104 4870 5582 4922
rect 5634 4870 5646 4922
rect 5698 4870 5710 4922
rect 5762 4870 5774 4922
rect 5826 4870 5838 4922
rect 5890 4870 14846 4922
rect 14898 4870 14910 4922
rect 14962 4870 14974 4922
rect 15026 4870 15038 4922
rect 15090 4870 15102 4922
rect 15154 4870 24110 4922
rect 24162 4870 24174 4922
rect 24226 4870 24238 4922
rect 24290 4870 24302 4922
rect 24354 4870 24366 4922
rect 24418 4870 28888 4922
rect 1104 4848 28888 4870
rect 9861 4811 9919 4817
rect 9861 4777 9873 4811
rect 9907 4808 9919 4811
rect 10134 4808 10140 4820
rect 9907 4780 10140 4808
rect 9907 4777 9919 4780
rect 9861 4771 9919 4777
rect 10134 4768 10140 4780
rect 10192 4768 10198 4820
rect 12618 4768 12624 4820
rect 12676 4808 12682 4820
rect 12986 4808 12992 4820
rect 12676 4780 12992 4808
rect 12676 4768 12682 4780
rect 12986 4768 12992 4780
rect 13044 4808 13050 4820
rect 13173 4811 13231 4817
rect 13173 4808 13185 4811
rect 13044 4780 13185 4808
rect 13044 4768 13050 4780
rect 13173 4777 13185 4780
rect 13219 4777 13231 4811
rect 13173 4771 13231 4777
rect 16485 4811 16543 4817
rect 16485 4777 16497 4811
rect 16531 4808 16543 4811
rect 17402 4808 17408 4820
rect 16531 4780 17408 4808
rect 16531 4777 16543 4780
rect 16485 4771 16543 4777
rect 17402 4768 17408 4780
rect 17460 4768 17466 4820
rect 18138 4808 18144 4820
rect 18099 4780 18144 4808
rect 18138 4768 18144 4780
rect 18196 4768 18202 4820
rect 20349 4811 20407 4817
rect 20349 4777 20361 4811
rect 20395 4808 20407 4811
rect 20530 4808 20536 4820
rect 20395 4780 20536 4808
rect 20395 4777 20407 4780
rect 20349 4771 20407 4777
rect 20530 4768 20536 4780
rect 20588 4768 20594 4820
rect 20993 4811 21051 4817
rect 20993 4777 21005 4811
rect 21039 4808 21051 4811
rect 23106 4808 23112 4820
rect 21039 4780 23112 4808
rect 21039 4777 21051 4780
rect 20993 4771 21051 4777
rect 23106 4768 23112 4780
rect 23164 4768 23170 4820
rect 12250 4700 12256 4752
rect 12308 4740 12314 4752
rect 13354 4740 13360 4752
rect 12308 4712 13360 4740
rect 12308 4700 12314 4712
rect 13354 4700 13360 4712
rect 13412 4740 13418 4752
rect 15197 4743 15255 4749
rect 15197 4740 15209 4743
rect 13412 4712 15209 4740
rect 13412 4700 13418 4712
rect 15197 4709 15209 4712
rect 15243 4740 15255 4743
rect 22649 4743 22707 4749
rect 15243 4712 22094 4740
rect 15243 4709 15255 4712
rect 15197 4703 15255 4709
rect 10134 4672 10140 4684
rect 9692 4644 10140 4672
rect 9306 4564 9312 4616
rect 9364 4604 9370 4616
rect 9692 4613 9720 4644
rect 10134 4632 10140 4644
rect 10192 4672 10198 4684
rect 10192 4644 10640 4672
rect 10192 4632 10198 4644
rect 9677 4607 9735 4613
rect 9677 4604 9689 4607
rect 9364 4576 9689 4604
rect 9364 4564 9370 4576
rect 9677 4573 9689 4576
rect 9723 4573 9735 4607
rect 10410 4604 10416 4616
rect 10371 4576 10416 4604
rect 9677 4567 9735 4573
rect 10410 4564 10416 4576
rect 10468 4564 10474 4616
rect 10612 4613 10640 4644
rect 11606 4632 11612 4684
rect 11664 4672 11670 4684
rect 11664 4644 12756 4672
rect 11664 4632 11670 4644
rect 10597 4607 10655 4613
rect 10597 4573 10609 4607
rect 10643 4573 10655 4607
rect 10597 4567 10655 4573
rect 10778 4564 10784 4616
rect 10836 4604 10842 4616
rect 11057 4607 11115 4613
rect 11057 4604 11069 4607
rect 10836 4576 11069 4604
rect 10836 4564 10842 4576
rect 11057 4573 11069 4576
rect 11103 4573 11115 4607
rect 11422 4604 11428 4616
rect 11383 4576 11428 4604
rect 11057 4567 11115 4573
rect 11422 4564 11428 4576
rect 11480 4564 11486 4616
rect 12158 4564 12164 4616
rect 12216 4604 12222 4616
rect 12437 4607 12495 4613
rect 12437 4604 12449 4607
rect 12216 4576 12449 4604
rect 12216 4564 12222 4576
rect 12437 4573 12449 4576
rect 12483 4573 12495 4607
rect 12437 4567 12495 4573
rect 12618 4564 12624 4616
rect 12676 4564 12682 4616
rect 12728 4613 12756 4644
rect 12894 4632 12900 4684
rect 12952 4672 12958 4684
rect 13265 4675 13323 4681
rect 13265 4672 13277 4675
rect 12952 4644 13277 4672
rect 12952 4632 12958 4644
rect 13265 4641 13277 4644
rect 13311 4672 13323 4675
rect 14369 4675 14427 4681
rect 14369 4672 14381 4675
rect 13311 4644 14381 4672
rect 13311 4641 13323 4644
rect 13265 4635 13323 4641
rect 14369 4641 14381 4644
rect 14415 4641 14427 4675
rect 14369 4635 14427 4641
rect 14734 4632 14740 4684
rect 14792 4672 14798 4684
rect 21174 4672 21180 4684
rect 14792 4644 19380 4672
rect 14792 4632 14798 4644
rect 12713 4607 12771 4613
rect 12713 4573 12725 4607
rect 12759 4573 12771 4607
rect 13170 4604 13176 4616
rect 13131 4576 13176 4604
rect 12713 4567 12771 4573
rect 9493 4539 9551 4545
rect 9493 4505 9505 4539
rect 9539 4536 9551 4539
rect 10796 4536 10824 4564
rect 9539 4508 10824 4536
rect 11609 4539 11667 4545
rect 9539 4505 9551 4508
rect 9493 4499 9551 4505
rect 11609 4505 11621 4539
rect 11655 4536 11667 4539
rect 12636 4536 12664 4564
rect 11655 4508 12664 4536
rect 12728 4536 12756 4567
rect 13170 4564 13176 4576
rect 13228 4564 13234 4616
rect 14090 4604 14096 4616
rect 14051 4576 14096 4604
rect 14090 4564 14096 4576
rect 14148 4564 14154 4616
rect 14550 4564 14556 4616
rect 14608 4604 14614 4616
rect 15565 4607 15623 4613
rect 15565 4604 15577 4607
rect 14608 4576 15577 4604
rect 14608 4564 14614 4576
rect 15565 4573 15577 4576
rect 15611 4573 15623 4607
rect 16114 4604 16120 4616
rect 16075 4576 16120 4604
rect 15565 4567 15623 4573
rect 16114 4564 16120 4576
rect 16172 4564 16178 4616
rect 16485 4607 16543 4613
rect 16485 4573 16497 4607
rect 16531 4604 16543 4607
rect 17218 4604 17224 4616
rect 16531 4576 17224 4604
rect 16531 4573 16543 4576
rect 16485 4567 16543 4573
rect 17218 4564 17224 4576
rect 17276 4564 17282 4616
rect 18414 4604 18420 4616
rect 18375 4576 18420 4604
rect 18414 4564 18420 4576
rect 18472 4564 18478 4616
rect 18693 4607 18751 4613
rect 18693 4573 18705 4607
rect 18739 4604 18751 4607
rect 18966 4604 18972 4616
rect 18739 4576 18972 4604
rect 18739 4573 18751 4576
rect 18693 4567 18751 4573
rect 18966 4564 18972 4576
rect 19024 4564 19030 4616
rect 19352 4613 19380 4644
rect 19444 4644 21180 4672
rect 19444 4613 19472 4644
rect 21174 4632 21180 4644
rect 21232 4632 21238 4684
rect 21821 4675 21879 4681
rect 21821 4641 21833 4675
rect 21867 4672 21879 4675
rect 21910 4672 21916 4684
rect 21867 4644 21916 4672
rect 21867 4641 21879 4644
rect 21821 4635 21879 4641
rect 21910 4632 21916 4644
rect 21968 4632 21974 4684
rect 22066 4672 22094 4712
rect 22649 4709 22661 4743
rect 22695 4740 22707 4743
rect 23934 4740 23940 4752
rect 22695 4712 23940 4740
rect 22695 4709 22707 4712
rect 22649 4703 22707 4709
rect 23934 4700 23940 4712
rect 23992 4700 23998 4752
rect 23014 4672 23020 4684
rect 22066 4644 23020 4672
rect 23014 4632 23020 4644
rect 23072 4672 23078 4684
rect 23072 4644 23428 4672
rect 23072 4632 23078 4644
rect 19337 4607 19395 4613
rect 19337 4573 19349 4607
rect 19383 4573 19395 4607
rect 19337 4567 19395 4573
rect 19429 4607 19487 4613
rect 19429 4573 19441 4607
rect 19475 4573 19487 4607
rect 19429 4567 19487 4573
rect 19705 4607 19763 4613
rect 19705 4573 19717 4607
rect 19751 4573 19763 4607
rect 19705 4567 19763 4573
rect 19797 4607 19855 4613
rect 19797 4573 19809 4607
rect 19843 4604 19855 4607
rect 20346 4604 20352 4616
rect 19843 4576 20352 4604
rect 19843 4573 19855 4576
rect 19797 4567 19855 4573
rect 13449 4539 13507 4545
rect 13449 4536 13461 4539
rect 12728 4508 13461 4536
rect 11655 4505 11667 4508
rect 11609 4499 11667 4505
rect 13449 4505 13461 4508
rect 13495 4505 13507 4539
rect 13449 4499 13507 4505
rect 15286 4496 15292 4548
rect 15344 4536 15350 4548
rect 15381 4539 15439 4545
rect 15381 4536 15393 4539
rect 15344 4508 15393 4536
rect 15344 4496 15350 4508
rect 15381 4505 15393 4508
rect 15427 4505 15439 4539
rect 17770 4536 17776 4548
rect 17731 4508 17776 4536
rect 15381 4499 15439 4505
rect 17770 4496 17776 4508
rect 17828 4496 17834 4548
rect 17957 4539 18015 4545
rect 17957 4505 17969 4539
rect 18003 4536 18015 4539
rect 18138 4536 18144 4548
rect 18003 4508 18144 4536
rect 18003 4505 18015 4508
rect 17957 4499 18015 4505
rect 18138 4496 18144 4508
rect 18196 4496 18202 4548
rect 18782 4536 18788 4548
rect 18695 4508 18788 4536
rect 18782 4496 18788 4508
rect 18840 4536 18846 4548
rect 19444 4536 19472 4567
rect 18840 4508 19472 4536
rect 19521 4539 19579 4545
rect 18840 4496 18846 4508
rect 19521 4505 19533 4539
rect 19567 4505 19579 4539
rect 19720 4536 19748 4567
rect 20346 4564 20352 4576
rect 20404 4564 20410 4616
rect 20530 4564 20536 4616
rect 20588 4604 20594 4616
rect 20809 4607 20867 4613
rect 20809 4604 20821 4607
rect 20588 4576 20821 4604
rect 20588 4564 20594 4576
rect 20809 4573 20821 4576
rect 20855 4573 20867 4607
rect 20809 4567 20867 4573
rect 21085 4607 21143 4613
rect 21085 4573 21097 4607
rect 21131 4604 21143 4607
rect 21361 4607 21419 4613
rect 21361 4604 21373 4607
rect 21131 4576 21373 4604
rect 21131 4573 21143 4576
rect 21085 4567 21143 4573
rect 21361 4573 21373 4576
rect 21407 4573 21419 4607
rect 21542 4604 21548 4616
rect 21503 4576 21548 4604
rect 21361 4567 21419 4573
rect 21542 4564 21548 4576
rect 21600 4564 21606 4616
rect 21729 4607 21787 4613
rect 21729 4573 21741 4607
rect 21775 4573 21787 4607
rect 21729 4567 21787 4573
rect 19978 4536 19984 4548
rect 19720 4508 19984 4536
rect 19521 4499 19579 4505
rect 12618 4428 12624 4480
rect 12676 4468 12682 4480
rect 12989 4471 13047 4477
rect 12989 4468 13001 4471
rect 12676 4440 13001 4468
rect 12676 4428 12682 4440
rect 12989 4437 13001 4440
rect 13035 4437 13047 4471
rect 16666 4468 16672 4480
rect 16627 4440 16672 4468
rect 12989 4431 13047 4437
rect 16666 4428 16672 4440
rect 16724 4428 16730 4480
rect 19334 4428 19340 4480
rect 19392 4468 19398 4480
rect 19536 4468 19564 4499
rect 19978 4496 19984 4508
rect 20036 4496 20042 4548
rect 21744 4536 21772 4567
rect 22554 4564 22560 4616
rect 22612 4604 22618 4616
rect 22649 4607 22707 4613
rect 22649 4604 22661 4607
rect 22612 4576 22661 4604
rect 22612 4564 22618 4576
rect 22649 4573 22661 4576
rect 22695 4573 22707 4607
rect 22649 4567 22707 4573
rect 22738 4564 22744 4616
rect 22796 4604 22802 4616
rect 23293 4607 23351 4613
rect 23293 4604 23305 4607
rect 22796 4576 22841 4604
rect 22940 4576 23305 4604
rect 22796 4564 22802 4576
rect 21818 4536 21824 4548
rect 21744 4508 21824 4536
rect 21818 4496 21824 4508
rect 21876 4496 21882 4548
rect 22002 4496 22008 4548
rect 22060 4536 22066 4548
rect 22940 4536 22968 4576
rect 23293 4573 23305 4576
rect 23339 4573 23351 4607
rect 23293 4567 23351 4573
rect 22060 4508 22968 4536
rect 23017 4539 23075 4545
rect 22060 4496 22066 4508
rect 23017 4505 23029 4539
rect 23063 4536 23075 4539
rect 23400 4536 23428 4644
rect 28350 4604 28356 4616
rect 28311 4576 28356 4604
rect 28350 4564 28356 4576
rect 28408 4564 28414 4616
rect 23063 4508 23428 4536
rect 23063 4505 23075 4508
rect 23017 4499 23075 4505
rect 19392 4440 19564 4468
rect 19797 4471 19855 4477
rect 19392 4428 19398 4440
rect 19797 4437 19809 4471
rect 19843 4468 19855 4471
rect 20070 4468 20076 4480
rect 19843 4440 20076 4468
rect 19843 4437 19855 4440
rect 19797 4431 19855 4437
rect 20070 4428 20076 4440
rect 20128 4428 20134 4480
rect 20622 4468 20628 4480
rect 20583 4440 20628 4468
rect 20622 4428 20628 4440
rect 20680 4428 20686 4480
rect 22925 4471 22983 4477
rect 22925 4437 22937 4471
rect 22971 4468 22983 4471
rect 23385 4471 23443 4477
rect 23385 4468 23397 4471
rect 22971 4440 23397 4468
rect 22971 4437 22983 4440
rect 22925 4431 22983 4437
rect 23385 4437 23397 4440
rect 23431 4437 23443 4471
rect 23385 4431 23443 4437
rect 1104 4378 28888 4400
rect 1104 4326 10214 4378
rect 10266 4326 10278 4378
rect 10330 4326 10342 4378
rect 10394 4326 10406 4378
rect 10458 4326 10470 4378
rect 10522 4326 19478 4378
rect 19530 4326 19542 4378
rect 19594 4326 19606 4378
rect 19658 4326 19670 4378
rect 19722 4326 19734 4378
rect 19786 4326 28888 4378
rect 1104 4304 28888 4326
rect 9769 4267 9827 4273
rect 9769 4233 9781 4267
rect 9815 4264 9827 4267
rect 9815 4236 10456 4264
rect 9815 4233 9827 4236
rect 9769 4227 9827 4233
rect 8110 4088 8116 4140
rect 8168 4128 8174 4140
rect 8389 4131 8447 4137
rect 8389 4128 8401 4131
rect 8168 4100 8401 4128
rect 8168 4088 8174 4100
rect 8389 4097 8401 4100
rect 8435 4097 8447 4131
rect 8389 4091 8447 4097
rect 8656 4131 8714 4137
rect 8656 4097 8668 4131
rect 8702 4128 8714 4131
rect 9950 4128 9956 4140
rect 8702 4100 9956 4128
rect 8702 4097 8714 4100
rect 8656 4091 8714 4097
rect 9950 4088 9956 4100
rect 10008 4088 10014 4140
rect 10428 4137 10456 4236
rect 11698 4224 11704 4276
rect 11756 4264 11762 4276
rect 12802 4264 12808 4276
rect 11756 4236 12808 4264
rect 11756 4224 11762 4236
rect 10229 4131 10287 4137
rect 10229 4097 10241 4131
rect 10275 4097 10287 4131
rect 10229 4091 10287 4097
rect 10413 4131 10471 4137
rect 10413 4097 10425 4131
rect 10459 4128 10471 4131
rect 10594 4128 10600 4140
rect 10459 4100 10600 4128
rect 10459 4097 10471 4100
rect 10413 4091 10471 4097
rect 10244 4060 10272 4091
rect 10594 4088 10600 4100
rect 10652 4088 10658 4140
rect 11793 4131 11851 4137
rect 11793 4097 11805 4131
rect 11839 4128 11851 4131
rect 12158 4128 12164 4140
rect 11839 4100 12164 4128
rect 11839 4097 11851 4100
rect 11793 4091 11851 4097
rect 12158 4088 12164 4100
rect 12216 4088 12222 4140
rect 12250 4088 12256 4140
rect 12308 4128 12314 4140
rect 12544 4137 12572 4236
rect 12802 4224 12808 4236
rect 12860 4224 12866 4276
rect 14001 4267 14059 4273
rect 14001 4264 14013 4267
rect 13648 4236 14013 4264
rect 13648 4205 13676 4236
rect 14001 4233 14013 4236
rect 14047 4264 14059 4267
rect 14090 4264 14096 4276
rect 14047 4236 14096 4264
rect 14047 4233 14059 4236
rect 14001 4227 14059 4233
rect 14090 4224 14096 4236
rect 14148 4224 14154 4276
rect 19334 4224 19340 4276
rect 19392 4264 19398 4276
rect 19429 4267 19487 4273
rect 19429 4264 19441 4267
rect 19392 4236 19441 4264
rect 19392 4224 19398 4236
rect 19429 4233 19441 4236
rect 19475 4233 19487 4267
rect 19429 4227 19487 4233
rect 21453 4267 21511 4273
rect 21453 4233 21465 4267
rect 21499 4264 21511 4267
rect 21542 4264 21548 4276
rect 21499 4236 21548 4264
rect 21499 4233 21511 4236
rect 21453 4227 21511 4233
rect 21542 4224 21548 4236
rect 21600 4224 21606 4276
rect 13633 4199 13691 4205
rect 13633 4165 13645 4199
rect 13679 4165 13691 4199
rect 13633 4159 13691 4165
rect 14182 4156 14188 4208
rect 14240 4196 14246 4208
rect 15114 4199 15172 4205
rect 15114 4196 15126 4199
rect 14240 4168 15126 4196
rect 14240 4156 14246 4168
rect 15114 4165 15126 4168
rect 15160 4165 15172 4199
rect 15114 4159 15172 4165
rect 16945 4199 17003 4205
rect 16945 4165 16957 4199
rect 16991 4196 17003 4199
rect 17034 4196 17040 4208
rect 16991 4168 17040 4196
rect 16991 4165 17003 4168
rect 16945 4159 17003 4165
rect 17034 4156 17040 4168
rect 17092 4156 17098 4208
rect 18966 4196 18972 4208
rect 17236 4168 17908 4196
rect 18927 4168 18972 4196
rect 17236 4140 17264 4168
rect 12391 4131 12449 4137
rect 12308 4100 12353 4128
rect 12308 4088 12314 4100
rect 12391 4097 12403 4131
rect 12437 4097 12449 4131
rect 12391 4091 12449 4097
rect 12529 4131 12587 4137
rect 12529 4097 12541 4131
rect 12575 4097 12587 4131
rect 12529 4091 12587 4097
rect 10778 4060 10784 4072
rect 10244 4032 10784 4060
rect 10778 4020 10784 4032
rect 10836 4020 10842 4072
rect 11701 4063 11759 4069
rect 11701 4029 11713 4063
rect 11747 4060 11759 4063
rect 12406 4060 12434 4091
rect 12618 4088 12624 4140
rect 12676 4128 12682 4140
rect 12676 4100 12721 4128
rect 12676 4088 12682 4100
rect 12894 4088 12900 4140
rect 12952 4128 12958 4140
rect 13170 4128 13176 4140
rect 12952 4100 13176 4128
rect 12952 4088 12958 4100
rect 13170 4088 13176 4100
rect 13228 4128 13234 4140
rect 13357 4131 13415 4137
rect 13357 4128 13369 4131
rect 13228 4100 13369 4128
rect 13228 4088 13234 4100
rect 13357 4097 13369 4100
rect 13403 4097 13415 4131
rect 16666 4128 16672 4140
rect 16627 4100 16672 4128
rect 13357 4091 13415 4097
rect 16666 4088 16672 4100
rect 16724 4088 16730 4140
rect 16761 4131 16819 4137
rect 16761 4097 16773 4131
rect 16807 4097 16819 4131
rect 17218 4128 17224 4140
rect 17179 4100 17224 4128
rect 16761 4091 16819 4097
rect 11747 4032 12434 4060
rect 11747 4029 11759 4032
rect 11701 4023 11759 4029
rect 12986 4020 12992 4072
rect 13044 4060 13050 4072
rect 13449 4063 13507 4069
rect 13449 4060 13461 4063
rect 13044 4032 13461 4060
rect 13044 4020 13050 4032
rect 13449 4029 13461 4032
rect 13495 4029 13507 4063
rect 15378 4060 15384 4072
rect 15339 4032 15384 4060
rect 13449 4023 13507 4029
rect 15378 4020 15384 4032
rect 15436 4020 15442 4072
rect 16776 4060 16804 4091
rect 17218 4088 17224 4100
rect 17276 4088 17282 4140
rect 17402 4128 17408 4140
rect 17363 4100 17408 4128
rect 17402 4088 17408 4100
rect 17460 4088 17466 4140
rect 17681 4131 17739 4137
rect 17681 4097 17693 4131
rect 17727 4128 17739 4131
rect 17770 4128 17776 4140
rect 17727 4100 17776 4128
rect 17727 4097 17739 4100
rect 17681 4091 17739 4097
rect 17770 4088 17776 4100
rect 17828 4088 17834 4140
rect 17880 4128 17908 4168
rect 18966 4156 18972 4168
rect 19024 4156 19030 4208
rect 20340 4199 20398 4205
rect 20340 4165 20352 4199
rect 20386 4196 20398 4199
rect 20622 4196 20628 4208
rect 20386 4168 20628 4196
rect 20386 4165 20398 4168
rect 20340 4159 20398 4165
rect 20622 4156 20628 4168
rect 20680 4156 20686 4208
rect 21910 4156 21916 4208
rect 21968 4196 21974 4208
rect 21968 4168 22048 4196
rect 21968 4156 21974 4168
rect 17957 4131 18015 4137
rect 17957 4128 17969 4131
rect 17880 4100 17969 4128
rect 17957 4097 17969 4100
rect 18003 4097 18015 4131
rect 17957 4091 18015 4097
rect 17313 4063 17371 4069
rect 17313 4060 17325 4063
rect 16776 4032 17325 4060
rect 17313 4029 17325 4032
rect 17359 4029 17371 4063
rect 17313 4023 17371 4029
rect 11422 3952 11428 4004
rect 11480 3992 11486 4004
rect 13173 3995 13231 4001
rect 13173 3992 13185 3995
rect 11480 3964 13185 3992
rect 11480 3952 11486 3964
rect 13173 3961 13185 3964
rect 13219 3961 13231 3995
rect 13173 3955 13231 3961
rect 10134 3884 10140 3936
rect 10192 3924 10198 3936
rect 10229 3927 10287 3933
rect 10229 3924 10241 3927
rect 10192 3896 10241 3924
rect 10192 3884 10198 3896
rect 10229 3893 10241 3896
rect 10275 3893 10287 3927
rect 10229 3887 10287 3893
rect 10597 3927 10655 3933
rect 10597 3893 10609 3927
rect 10643 3924 10655 3927
rect 11606 3924 11612 3936
rect 10643 3896 11612 3924
rect 10643 3893 10655 3896
rect 10597 3887 10655 3893
rect 11606 3884 11612 3896
rect 11664 3884 11670 3936
rect 11790 3884 11796 3936
rect 11848 3924 11854 3936
rect 12069 3927 12127 3933
rect 12069 3924 12081 3927
rect 11848 3896 12081 3924
rect 11848 3884 11854 3896
rect 12069 3893 12081 3896
rect 12115 3893 12127 3927
rect 12069 3887 12127 3893
rect 12158 3884 12164 3936
rect 12216 3924 12222 3936
rect 12894 3924 12900 3936
rect 12216 3896 12900 3924
rect 12216 3884 12222 3896
rect 12894 3884 12900 3896
rect 12952 3884 12958 3936
rect 13262 3884 13268 3936
rect 13320 3924 13326 3936
rect 13357 3927 13415 3933
rect 13357 3924 13369 3927
rect 13320 3896 13369 3924
rect 13320 3884 13326 3896
rect 13357 3893 13369 3896
rect 13403 3893 13415 3927
rect 16942 3924 16948 3936
rect 16903 3896 16948 3924
rect 13357 3887 13415 3893
rect 16942 3884 16948 3896
rect 17000 3884 17006 3936
rect 17972 3924 18000 4091
rect 18138 4088 18144 4140
rect 18196 4128 18202 4140
rect 19245 4131 19303 4137
rect 19245 4128 19257 4131
rect 18196 4100 19257 4128
rect 18196 4088 18202 4100
rect 19245 4097 19257 4100
rect 19291 4128 19303 4131
rect 19702 4128 19708 4140
rect 19291 4100 19708 4128
rect 19291 4097 19303 4100
rect 19245 4091 19303 4097
rect 19702 4088 19708 4100
rect 19760 4088 19766 4140
rect 19886 4088 19892 4140
rect 19944 4128 19950 4140
rect 22020 4137 22048 4168
rect 20073 4131 20131 4137
rect 20073 4128 20085 4131
rect 19944 4100 20085 4128
rect 19944 4088 19950 4100
rect 20073 4097 20085 4100
rect 20119 4097 20131 4131
rect 20073 4091 20131 4097
rect 22005 4131 22063 4137
rect 22005 4097 22017 4131
rect 22051 4097 22063 4131
rect 22005 4091 22063 4097
rect 18598 4020 18604 4072
rect 18656 4060 18662 4072
rect 19061 4063 19119 4069
rect 19061 4060 19073 4063
rect 18656 4032 19073 4060
rect 18656 4020 18662 4032
rect 19061 4029 19073 4032
rect 19107 4029 19119 4063
rect 21910 4060 21916 4072
rect 21871 4032 21916 4060
rect 19061 4023 19119 4029
rect 21910 4020 21916 4032
rect 21968 4020 21974 4072
rect 22020 3992 22048 4091
rect 23934 4088 23940 4140
rect 23992 4137 23998 4140
rect 23992 4128 24004 4137
rect 23992 4100 24037 4128
rect 23992 4091 24004 4100
rect 23992 4088 23998 4091
rect 22373 4063 22431 4069
rect 22373 4029 22385 4063
rect 22419 4060 22431 4063
rect 22738 4060 22744 4072
rect 22419 4032 22744 4060
rect 22419 4029 22431 4032
rect 22373 4023 22431 4029
rect 22738 4020 22744 4032
rect 22796 4020 22802 4072
rect 24213 4063 24271 4069
rect 24213 4029 24225 4063
rect 24259 4060 24271 4063
rect 24486 4060 24492 4072
rect 24259 4032 24492 4060
rect 24259 4029 24271 4032
rect 24213 4023 24271 4029
rect 24486 4020 24492 4032
rect 24544 4020 24550 4072
rect 22833 3995 22891 4001
rect 22833 3992 22845 3995
rect 22020 3964 22845 3992
rect 22833 3961 22845 3964
rect 22879 3961 22891 3995
rect 22833 3955 22891 3961
rect 18969 3927 19027 3933
rect 18969 3924 18981 3927
rect 17972 3896 18981 3924
rect 18969 3893 18981 3896
rect 19015 3924 19027 3927
rect 19242 3924 19248 3936
rect 19015 3896 19248 3924
rect 19015 3893 19027 3896
rect 18969 3887 19027 3893
rect 19242 3884 19248 3896
rect 19300 3884 19306 3936
rect 1104 3834 28888 3856
rect 1104 3782 5582 3834
rect 5634 3782 5646 3834
rect 5698 3782 5710 3834
rect 5762 3782 5774 3834
rect 5826 3782 5838 3834
rect 5890 3782 14846 3834
rect 14898 3782 14910 3834
rect 14962 3782 14974 3834
rect 15026 3782 15038 3834
rect 15090 3782 15102 3834
rect 15154 3782 24110 3834
rect 24162 3782 24174 3834
rect 24226 3782 24238 3834
rect 24290 3782 24302 3834
rect 24354 3782 24366 3834
rect 24418 3782 28888 3834
rect 1104 3760 28888 3782
rect 11793 3723 11851 3729
rect 11793 3689 11805 3723
rect 11839 3720 11851 3723
rect 13078 3720 13084 3732
rect 11839 3692 13084 3720
rect 11839 3689 11851 3692
rect 11793 3683 11851 3689
rect 13078 3680 13084 3692
rect 13136 3680 13142 3732
rect 17589 3723 17647 3729
rect 17589 3689 17601 3723
rect 17635 3720 17647 3723
rect 17770 3720 17776 3732
rect 17635 3692 17776 3720
rect 17635 3689 17647 3692
rect 17589 3683 17647 3689
rect 17770 3680 17776 3692
rect 17828 3720 17834 3732
rect 17865 3723 17923 3729
rect 17865 3720 17877 3723
rect 17828 3692 17877 3720
rect 17828 3680 17834 3692
rect 17865 3689 17877 3692
rect 17911 3689 17923 3723
rect 17865 3683 17923 3689
rect 18325 3723 18383 3729
rect 18325 3689 18337 3723
rect 18371 3720 18383 3723
rect 18414 3720 18420 3732
rect 18371 3692 18420 3720
rect 18371 3689 18383 3692
rect 18325 3683 18383 3689
rect 18414 3680 18420 3692
rect 18472 3680 18478 3732
rect 18966 3680 18972 3732
rect 19024 3720 19030 3732
rect 19521 3723 19579 3729
rect 19521 3720 19533 3723
rect 19024 3692 19533 3720
rect 19024 3680 19030 3692
rect 19521 3689 19533 3692
rect 19567 3689 19579 3723
rect 19521 3683 19579 3689
rect 19981 3723 20039 3729
rect 19981 3689 19993 3723
rect 20027 3689 20039 3723
rect 19981 3683 20039 3689
rect 20349 3723 20407 3729
rect 20349 3689 20361 3723
rect 20395 3720 20407 3723
rect 21910 3720 21916 3732
rect 20395 3692 21916 3720
rect 20395 3689 20407 3692
rect 20349 3683 20407 3689
rect 12161 3655 12219 3661
rect 12161 3621 12173 3655
rect 12207 3652 12219 3655
rect 12250 3652 12256 3664
rect 12207 3624 12256 3652
rect 12207 3621 12219 3624
rect 12161 3615 12219 3621
rect 12250 3612 12256 3624
rect 12308 3612 12314 3664
rect 13262 3652 13268 3664
rect 12360 3624 13268 3652
rect 12360 3593 12388 3624
rect 13262 3612 13268 3624
rect 13320 3612 13326 3664
rect 13722 3652 13728 3664
rect 13683 3624 13728 3652
rect 13722 3612 13728 3624
rect 13780 3612 13786 3664
rect 19242 3612 19248 3664
rect 19300 3652 19306 3664
rect 19996 3652 20024 3683
rect 21910 3680 21916 3692
rect 21968 3680 21974 3732
rect 19300 3624 20024 3652
rect 19300 3612 19306 3624
rect 12345 3587 12403 3593
rect 10888 3556 12296 3584
rect 10888 3528 10916 3556
rect 10870 3516 10876 3528
rect 10831 3488 10876 3516
rect 10870 3476 10876 3488
rect 10928 3476 10934 3528
rect 11149 3519 11207 3525
rect 11149 3485 11161 3519
rect 11195 3516 11207 3519
rect 11790 3516 11796 3528
rect 11195 3488 11796 3516
rect 11195 3485 11207 3488
rect 11149 3479 11207 3485
rect 11790 3476 11796 3488
rect 11848 3476 11854 3528
rect 11882 3476 11888 3528
rect 11940 3516 11946 3528
rect 12069 3519 12127 3525
rect 12069 3516 12081 3519
rect 11940 3488 12081 3516
rect 11940 3476 11946 3488
rect 12069 3485 12081 3488
rect 12115 3485 12127 3519
rect 12268 3516 12296 3556
rect 12345 3553 12357 3587
rect 12391 3553 12403 3587
rect 12345 3547 12403 3553
rect 12434 3544 12440 3596
rect 12492 3584 12498 3596
rect 13170 3584 13176 3596
rect 12492 3556 13032 3584
rect 13131 3556 13176 3584
rect 12492 3544 12498 3556
rect 12268 3488 12572 3516
rect 12069 3479 12127 3485
rect 11422 3448 11428 3460
rect 11383 3420 11428 3448
rect 11422 3408 11428 3420
rect 11480 3408 11486 3460
rect 11606 3448 11612 3460
rect 11567 3420 11612 3448
rect 11606 3408 11612 3420
rect 11664 3408 11670 3460
rect 12345 3451 12403 3457
rect 12345 3448 12357 3451
rect 11716 3420 12357 3448
rect 10962 3380 10968 3392
rect 11020 3389 11026 3392
rect 10929 3352 10968 3380
rect 10962 3340 10968 3352
rect 11020 3343 11029 3389
rect 11057 3383 11115 3389
rect 11057 3349 11069 3383
rect 11103 3380 11115 3383
rect 11716 3380 11744 3420
rect 12345 3417 12357 3420
rect 12391 3417 12403 3451
rect 12544 3448 12572 3488
rect 12618 3476 12624 3528
rect 12676 3516 12682 3528
rect 13004 3525 13032 3556
rect 13170 3544 13176 3556
rect 13228 3544 13234 3596
rect 13538 3584 13544 3596
rect 13280 3556 13544 3584
rect 12897 3519 12955 3525
rect 12897 3516 12909 3519
rect 12676 3488 12909 3516
rect 12676 3476 12682 3488
rect 12897 3485 12909 3488
rect 12943 3485 12955 3519
rect 12897 3479 12955 3485
rect 12989 3519 13047 3525
rect 12989 3485 13001 3519
rect 13035 3516 13047 3519
rect 13280 3516 13308 3556
rect 13538 3544 13544 3556
rect 13596 3544 13602 3596
rect 18049 3587 18107 3593
rect 18049 3553 18061 3587
rect 18095 3584 18107 3587
rect 18598 3584 18604 3596
rect 18095 3556 18604 3584
rect 18095 3553 18107 3556
rect 18049 3547 18107 3553
rect 18598 3544 18604 3556
rect 18656 3584 18662 3596
rect 19383 3587 19441 3593
rect 19383 3584 19395 3587
rect 18656 3556 19395 3584
rect 18656 3544 18662 3556
rect 19383 3553 19395 3556
rect 19429 3553 19441 3587
rect 19383 3547 19441 3553
rect 19536 3556 19840 3584
rect 13446 3516 13452 3528
rect 13035 3488 13308 3516
rect 13407 3488 13452 3516
rect 13035 3485 13047 3488
rect 12989 3479 13047 3485
rect 13446 3476 13452 3488
rect 13504 3476 13510 3528
rect 16209 3519 16267 3525
rect 16209 3485 16221 3519
rect 16255 3516 16267 3519
rect 16758 3516 16764 3528
rect 16255 3488 16764 3516
rect 16255 3485 16267 3488
rect 16209 3479 16267 3485
rect 16758 3476 16764 3488
rect 16816 3476 16822 3528
rect 17865 3519 17923 3525
rect 17865 3485 17877 3519
rect 17911 3516 17923 3519
rect 17954 3516 17960 3528
rect 17911 3488 17960 3516
rect 17911 3485 17923 3488
rect 17865 3479 17923 3485
rect 17954 3476 17960 3488
rect 18012 3476 18018 3528
rect 18138 3516 18144 3528
rect 18099 3488 18144 3516
rect 18138 3476 18144 3488
rect 18196 3476 18202 3528
rect 19242 3516 19248 3528
rect 19203 3488 19248 3516
rect 19242 3476 19248 3488
rect 19300 3476 19306 3528
rect 13725 3451 13783 3457
rect 13725 3448 13737 3451
rect 12544 3420 13737 3448
rect 12345 3411 12403 3417
rect 13725 3417 13737 3420
rect 13771 3448 13783 3451
rect 13998 3448 14004 3460
rect 13771 3420 14004 3448
rect 13771 3417 13783 3420
rect 13725 3411 13783 3417
rect 13998 3408 14004 3420
rect 14056 3408 14062 3460
rect 16476 3451 16534 3457
rect 16476 3417 16488 3451
rect 16522 3448 16534 3451
rect 16942 3448 16948 3460
rect 16522 3420 16948 3448
rect 16522 3417 16534 3420
rect 16476 3411 16534 3417
rect 16942 3408 16948 3420
rect 17000 3408 17006 3460
rect 11103 3352 11744 3380
rect 13173 3383 13231 3389
rect 11103 3349 11115 3352
rect 11057 3343 11115 3349
rect 13173 3349 13185 3383
rect 13219 3380 13231 3383
rect 13541 3383 13599 3389
rect 13541 3380 13553 3383
rect 13219 3352 13553 3380
rect 13219 3349 13231 3352
rect 13173 3343 13231 3349
rect 13541 3349 13553 3352
rect 13587 3349 13599 3383
rect 13541 3343 13599 3349
rect 11020 3340 11026 3343
rect 17402 3340 17408 3392
rect 17460 3380 17466 3392
rect 19536 3380 19564 3556
rect 19702 3516 19708 3528
rect 19663 3488 19708 3516
rect 19702 3476 19708 3488
rect 19760 3476 19766 3528
rect 19812 3516 19840 3556
rect 19886 3544 19892 3596
rect 19944 3584 19950 3596
rect 20717 3587 20775 3593
rect 20717 3584 20729 3587
rect 19944 3556 20729 3584
rect 19944 3544 19950 3556
rect 20717 3553 20729 3556
rect 20763 3553 20775 3587
rect 20717 3547 20775 3553
rect 19981 3519 20039 3525
rect 19981 3516 19993 3519
rect 19812 3488 19993 3516
rect 19981 3485 19993 3488
rect 20027 3485 20039 3519
rect 19981 3479 20039 3485
rect 20073 3519 20131 3525
rect 20073 3485 20085 3519
rect 20119 3485 20131 3519
rect 20073 3479 20131 3485
rect 20984 3519 21042 3525
rect 20984 3485 20996 3519
rect 21030 3516 21042 3519
rect 21450 3516 21456 3528
rect 21030 3488 21456 3516
rect 21030 3485 21042 3488
rect 20984 3479 21042 3485
rect 19720 3448 19748 3476
rect 20088 3448 20116 3479
rect 21450 3476 21456 3488
rect 21508 3476 21514 3528
rect 24397 3519 24455 3525
rect 24397 3485 24409 3519
rect 24443 3516 24455 3519
rect 24486 3516 24492 3528
rect 24443 3488 24492 3516
rect 24443 3485 24455 3488
rect 24397 3479 24455 3485
rect 24486 3476 24492 3488
rect 24544 3476 24550 3528
rect 20346 3448 20352 3460
rect 19720 3420 20352 3448
rect 20346 3408 20352 3420
rect 20404 3408 20410 3460
rect 22830 3408 22836 3460
rect 22888 3448 22894 3460
rect 24642 3451 24700 3457
rect 24642 3448 24654 3451
rect 22888 3420 24654 3448
rect 22888 3408 22894 3420
rect 24642 3417 24654 3420
rect 24688 3417 24700 3451
rect 24642 3411 24700 3417
rect 17460 3352 19564 3380
rect 19705 3383 19763 3389
rect 17460 3340 17466 3352
rect 19705 3349 19717 3383
rect 19751 3380 19763 3383
rect 19978 3380 19984 3392
rect 19751 3352 19984 3380
rect 19751 3349 19763 3352
rect 19705 3343 19763 3349
rect 19978 3340 19984 3352
rect 20036 3340 20042 3392
rect 22097 3383 22155 3389
rect 22097 3349 22109 3383
rect 22143 3380 22155 3383
rect 22278 3380 22284 3392
rect 22143 3352 22284 3380
rect 22143 3349 22155 3352
rect 22097 3343 22155 3349
rect 22278 3340 22284 3352
rect 22336 3340 22342 3392
rect 25777 3383 25835 3389
rect 25777 3349 25789 3383
rect 25823 3380 25835 3383
rect 28074 3380 28080 3392
rect 25823 3352 28080 3380
rect 25823 3349 25835 3352
rect 25777 3343 25835 3349
rect 28074 3340 28080 3352
rect 28132 3340 28138 3392
rect 1104 3290 28888 3312
rect 1104 3238 10214 3290
rect 10266 3238 10278 3290
rect 10330 3238 10342 3290
rect 10394 3238 10406 3290
rect 10458 3238 10470 3290
rect 10522 3238 19478 3290
rect 19530 3238 19542 3290
rect 19594 3238 19606 3290
rect 19658 3238 19670 3290
rect 19722 3238 19734 3290
rect 19786 3238 28888 3290
rect 1104 3216 28888 3238
rect 8202 3176 8208 3188
rect 8163 3148 8208 3176
rect 8202 3136 8208 3148
rect 8260 3136 8266 3188
rect 11974 3136 11980 3188
rect 12032 3136 12038 3188
rect 13170 3136 13176 3188
rect 13228 3176 13234 3188
rect 13357 3179 13415 3185
rect 13357 3176 13369 3179
rect 13228 3148 13369 3176
rect 13228 3136 13234 3148
rect 13357 3145 13369 3148
rect 13403 3145 13415 3179
rect 20346 3176 20352 3188
rect 20307 3148 20352 3176
rect 13357 3139 13415 3145
rect 20346 3136 20352 3148
rect 20404 3136 20410 3188
rect 7592 3111 7650 3117
rect 7592 3077 7604 3111
rect 7638 3108 7650 3111
rect 8220 3108 8248 3136
rect 11992 3108 12020 3136
rect 15378 3108 15384 3120
rect 7638 3080 8248 3108
rect 11716 3080 15384 3108
rect 7638 3077 7650 3080
rect 7592 3071 7650 3077
rect 7837 3043 7895 3049
rect 7837 3009 7849 3043
rect 7883 3040 7895 3043
rect 8110 3040 8116 3052
rect 7883 3012 8116 3040
rect 7883 3009 7895 3012
rect 7837 3003 7895 3009
rect 8110 3000 8116 3012
rect 8168 3000 8174 3052
rect 11716 3049 11744 3080
rect 11701 3043 11759 3049
rect 11701 3009 11713 3043
rect 11747 3009 11759 3043
rect 11957 3043 12015 3049
rect 11957 3040 11969 3043
rect 11701 3003 11759 3009
rect 11808 3012 11969 3040
rect 10962 2932 10968 2984
rect 11020 2972 11026 2984
rect 11808 2972 11836 3012
rect 11957 3009 11969 3012
rect 12003 3009 12015 3043
rect 11957 3003 12015 3009
rect 13722 3000 13728 3052
rect 13780 3040 13786 3052
rect 14752 3049 14780 3080
rect 15378 3068 15384 3080
rect 15436 3068 15442 3120
rect 19886 3108 19892 3120
rect 18984 3080 19892 3108
rect 18984 3049 19012 3080
rect 19886 3068 19892 3080
rect 19944 3068 19950 3120
rect 14470 3043 14528 3049
rect 14470 3040 14482 3043
rect 13780 3012 14482 3040
rect 13780 3000 13786 3012
rect 14470 3009 14482 3012
rect 14516 3009 14528 3043
rect 14470 3003 14528 3009
rect 14737 3043 14795 3049
rect 14737 3009 14749 3043
rect 14783 3009 14795 3043
rect 14737 3003 14795 3009
rect 18969 3043 19027 3049
rect 18969 3009 18981 3043
rect 19015 3009 19027 3043
rect 18969 3003 19027 3009
rect 19236 3043 19294 3049
rect 19236 3009 19248 3043
rect 19282 3040 19294 3043
rect 20070 3040 20076 3052
rect 19282 3012 20076 3040
rect 19282 3009 19294 3012
rect 19236 3003 19294 3009
rect 20070 3000 20076 3012
rect 20128 3000 20134 3052
rect 28074 3040 28080 3052
rect 28035 3012 28080 3040
rect 28074 3000 28080 3012
rect 28132 3000 28138 3052
rect 11020 2944 11836 2972
rect 11020 2932 11026 2944
rect 13081 2907 13139 2913
rect 13081 2873 13093 2907
rect 13127 2904 13139 2907
rect 13262 2904 13268 2916
rect 13127 2876 13268 2904
rect 13127 2873 13139 2876
rect 13081 2867 13139 2873
rect 13262 2864 13268 2876
rect 13320 2864 13326 2916
rect 1489 2839 1547 2845
rect 1489 2805 1501 2839
rect 1535 2836 1547 2839
rect 1670 2836 1676 2848
rect 1535 2808 1676 2836
rect 1535 2805 1547 2808
rect 1489 2799 1547 2805
rect 1670 2796 1676 2808
rect 1728 2796 1734 2848
rect 5902 2796 5908 2848
rect 5960 2836 5966 2848
rect 6457 2839 6515 2845
rect 6457 2836 6469 2839
rect 5960 2808 6469 2836
rect 5960 2796 5966 2808
rect 6457 2805 6469 2808
rect 6503 2805 6515 2839
rect 28258 2836 28264 2848
rect 28219 2808 28264 2836
rect 6457 2799 6515 2805
rect 28258 2796 28264 2808
rect 28316 2796 28322 2848
rect 1104 2746 28888 2768
rect 1104 2694 5582 2746
rect 5634 2694 5646 2746
rect 5698 2694 5710 2746
rect 5762 2694 5774 2746
rect 5826 2694 5838 2746
rect 5890 2694 14846 2746
rect 14898 2694 14910 2746
rect 14962 2694 14974 2746
rect 15026 2694 15038 2746
rect 15090 2694 15102 2746
rect 15154 2694 24110 2746
rect 24162 2694 24174 2746
rect 24226 2694 24238 2746
rect 24290 2694 24302 2746
rect 24354 2694 24366 2746
rect 24418 2694 28888 2746
rect 1104 2672 28888 2694
rect 17034 2632 17040 2644
rect 16995 2604 17040 2632
rect 17034 2592 17040 2604
rect 17092 2592 17098 2644
rect 20714 2632 20720 2644
rect 20675 2604 20720 2632
rect 20714 2592 20720 2604
rect 20772 2592 20778 2644
rect 1857 2567 1915 2573
rect 1857 2533 1869 2567
rect 1903 2564 1915 2567
rect 1903 2536 6914 2564
rect 1903 2533 1915 2536
rect 1857 2527 1915 2533
rect 5902 2496 5908 2508
rect 2424 2468 5908 2496
rect 2424 2437 2452 2468
rect 5902 2456 5908 2468
rect 5960 2456 5966 2508
rect 6886 2496 6914 2536
rect 20438 2524 20444 2576
rect 20496 2564 20502 2576
rect 27801 2567 27859 2573
rect 27801 2564 27813 2567
rect 20496 2536 27813 2564
rect 20496 2524 20502 2536
rect 27801 2533 27813 2536
rect 27847 2533 27859 2567
rect 27801 2527 27859 2533
rect 18506 2496 18512 2508
rect 6886 2468 18512 2496
rect 18506 2456 18512 2468
rect 18564 2456 18570 2508
rect 19521 2499 19579 2505
rect 19521 2465 19533 2499
rect 19567 2496 19579 2499
rect 20346 2496 20352 2508
rect 19567 2468 20352 2496
rect 19567 2465 19579 2468
rect 19521 2459 19579 2465
rect 20346 2456 20352 2468
rect 20404 2456 20410 2508
rect 2409 2431 2467 2437
rect 2409 2397 2421 2431
rect 2455 2397 2467 2431
rect 2409 2391 2467 2397
rect 3234 2388 3240 2440
rect 3292 2428 3298 2440
rect 3789 2431 3847 2437
rect 3789 2428 3801 2431
rect 3292 2400 3801 2428
rect 3292 2388 3298 2400
rect 3789 2397 3801 2400
rect 3835 2397 3847 2431
rect 3789 2391 3847 2397
rect 6454 2388 6460 2440
rect 6512 2428 6518 2440
rect 6549 2431 6607 2437
rect 6549 2428 6561 2431
rect 6512 2400 6561 2428
rect 6512 2388 6518 2400
rect 6549 2397 6561 2400
rect 6595 2397 6607 2431
rect 6549 2391 6607 2397
rect 12250 2388 12256 2440
rect 12308 2428 12314 2440
rect 12345 2431 12403 2437
rect 12345 2428 12357 2431
rect 12308 2400 12357 2428
rect 12308 2388 12314 2400
rect 12345 2397 12357 2400
rect 12391 2397 12403 2431
rect 19245 2431 19303 2437
rect 19245 2428 19257 2431
rect 12345 2391 12403 2397
rect 18800 2400 19257 2428
rect 1670 2360 1676 2372
rect 1631 2332 1676 2360
rect 1670 2320 1676 2332
rect 1728 2320 1734 2372
rect 5353 2363 5411 2369
rect 5353 2360 5365 2363
rect 5184 2332 5365 2360
rect 5184 2304 5212 2332
rect 5353 2329 5365 2332
rect 5399 2329 5411 2363
rect 5353 2323 5411 2329
rect 5721 2363 5779 2369
rect 5721 2329 5733 2363
rect 5767 2360 5779 2363
rect 15654 2360 15660 2372
rect 5767 2332 15660 2360
rect 5767 2329 5779 2332
rect 5721 2323 5779 2329
rect 15654 2320 15660 2332
rect 15712 2320 15718 2372
rect 16301 2363 16359 2369
rect 16301 2329 16313 2363
rect 16347 2360 16359 2363
rect 16758 2360 16764 2372
rect 16347 2332 16764 2360
rect 16347 2329 16359 2332
rect 16301 2323 16359 2329
rect 16758 2320 16764 2332
rect 16816 2360 16822 2372
rect 16945 2363 17003 2369
rect 16945 2360 16957 2363
rect 16816 2332 16957 2360
rect 16816 2320 16822 2332
rect 16945 2329 16957 2332
rect 16991 2329 17003 2363
rect 16945 2323 17003 2329
rect 2222 2292 2228 2304
rect 2183 2264 2228 2292
rect 2222 2252 2228 2264
rect 2280 2252 2286 2304
rect 4985 2295 5043 2301
rect 4985 2261 4997 2295
rect 5031 2292 5043 2295
rect 5166 2292 5172 2304
rect 5031 2264 5172 2292
rect 5031 2261 5043 2264
rect 4985 2255 5043 2261
rect 5166 2252 5172 2264
rect 5224 2252 5230 2304
rect 18690 2252 18696 2304
rect 18748 2292 18754 2304
rect 18800 2301 18828 2400
rect 19245 2397 19257 2400
rect 19291 2397 19303 2431
rect 19245 2391 19303 2397
rect 20714 2388 20720 2440
rect 20772 2428 20778 2440
rect 20901 2431 20959 2437
rect 20901 2428 20913 2431
rect 20772 2400 20913 2428
rect 20772 2388 20778 2400
rect 20901 2397 20913 2400
rect 20947 2428 20959 2431
rect 21177 2431 21235 2437
rect 21177 2428 21189 2431
rect 20947 2400 21189 2428
rect 20947 2397 20959 2400
rect 20901 2391 20959 2397
rect 21177 2397 21189 2400
rect 21223 2397 21235 2431
rect 22278 2428 22284 2440
rect 22239 2400 22284 2428
rect 21177 2391 21235 2397
rect 22278 2388 22284 2400
rect 22336 2388 22342 2440
rect 25222 2428 25228 2440
rect 25183 2400 25228 2428
rect 25222 2388 25228 2400
rect 25280 2388 25286 2440
rect 26418 2388 26424 2440
rect 26476 2428 26482 2440
rect 26973 2431 27031 2437
rect 26973 2428 26985 2431
rect 26476 2400 26985 2428
rect 26476 2388 26482 2400
rect 26973 2397 26985 2400
rect 27019 2397 27031 2431
rect 26973 2391 27031 2397
rect 27985 2363 28043 2369
rect 27985 2329 27997 2363
rect 28031 2329 28043 2363
rect 27985 2323 28043 2329
rect 18785 2295 18843 2301
rect 18785 2292 18797 2295
rect 18748 2264 18797 2292
rect 18748 2252 18754 2264
rect 18785 2261 18797 2264
rect 18831 2261 18843 2295
rect 18785 2255 18843 2261
rect 21910 2252 21916 2304
rect 21968 2292 21974 2304
rect 22097 2295 22155 2301
rect 22097 2292 22109 2295
rect 21968 2264 22109 2292
rect 21968 2252 21974 2264
rect 22097 2261 22109 2264
rect 22143 2261 22155 2295
rect 22097 2255 22155 2261
rect 25130 2252 25136 2304
rect 25188 2292 25194 2304
rect 25409 2295 25467 2301
rect 25409 2292 25421 2295
rect 25188 2264 25421 2292
rect 25188 2252 25194 2264
rect 25409 2261 25421 2264
rect 25455 2261 25467 2295
rect 25409 2255 25467 2261
rect 27525 2295 27583 2301
rect 27525 2261 27537 2295
rect 27571 2292 27583 2295
rect 27706 2292 27712 2304
rect 27571 2264 27712 2292
rect 27571 2261 27583 2264
rect 27525 2255 27583 2261
rect 27706 2252 27712 2264
rect 27764 2292 27770 2304
rect 28000 2292 28028 2323
rect 27764 2264 28028 2292
rect 27764 2252 27770 2264
rect 1104 2202 28888 2224
rect 1104 2150 10214 2202
rect 10266 2150 10278 2202
rect 10330 2150 10342 2202
rect 10394 2150 10406 2202
rect 10458 2150 10470 2202
rect 10522 2150 19478 2202
rect 19530 2150 19542 2202
rect 19594 2150 19606 2202
rect 19658 2150 19670 2202
rect 19722 2150 19734 2202
rect 19786 2150 28888 2202
rect 1104 2128 28888 2150
<< via1 >>
rect 5582 27718 5634 27770
rect 5646 27718 5698 27770
rect 5710 27718 5762 27770
rect 5774 27718 5826 27770
rect 5838 27718 5890 27770
rect 14846 27718 14898 27770
rect 14910 27718 14962 27770
rect 14974 27718 15026 27770
rect 15038 27718 15090 27770
rect 15102 27718 15154 27770
rect 24110 27718 24162 27770
rect 24174 27718 24226 27770
rect 24238 27718 24290 27770
rect 24302 27718 24354 27770
rect 24366 27718 24418 27770
rect 2412 27591 2464 27600
rect 2412 27557 2421 27591
rect 2421 27557 2455 27591
rect 2455 27557 2464 27591
rect 2412 27548 2464 27557
rect 3976 27591 4028 27600
rect 3976 27557 3985 27591
rect 3985 27557 4019 27591
rect 4019 27557 4028 27591
rect 3976 27548 4028 27557
rect 16488 27548 16540 27600
rect 19432 27591 19484 27600
rect 19432 27557 19441 27591
rect 19441 27557 19475 27591
rect 19475 27557 19484 27591
rect 19432 27548 19484 27557
rect 21272 27548 21324 27600
rect 22376 27591 22428 27600
rect 22376 27557 22385 27591
rect 22385 27557 22419 27591
rect 22419 27557 22428 27591
rect 22376 27548 22428 27557
rect 23940 27591 23992 27600
rect 23940 27557 23949 27591
rect 23949 27557 23983 27591
rect 23983 27557 23992 27591
rect 23940 27548 23992 27557
rect 25504 27591 25556 27600
rect 25504 27557 25513 27591
rect 25513 27557 25547 27591
rect 25547 27557 25556 27591
rect 25504 27548 25556 27557
rect 25872 27591 25924 27600
rect 25872 27557 25881 27591
rect 25881 27557 25915 27591
rect 25915 27557 25924 27591
rect 25872 27548 25924 27557
rect 27988 27548 28040 27600
rect 28264 27591 28316 27600
rect 28264 27557 28273 27591
rect 28273 27557 28307 27591
rect 28307 27557 28316 27591
rect 28264 27548 28316 27557
rect 1676 27455 1728 27464
rect 1676 27421 1685 27455
rect 1685 27421 1719 27455
rect 1719 27421 1728 27455
rect 1676 27412 1728 27421
rect 10508 27455 10560 27464
rect 10508 27421 10517 27455
rect 10517 27421 10551 27455
rect 10551 27421 10560 27455
rect 10508 27412 10560 27421
rect 18328 27412 18380 27464
rect 25136 27412 25188 27464
rect 3148 27387 3200 27396
rect 3148 27353 3157 27387
rect 3157 27353 3191 27387
rect 3191 27353 3200 27387
rect 3148 27344 3200 27353
rect 10784 27344 10836 27396
rect 25044 27387 25096 27396
rect 25044 27353 25053 27387
rect 25053 27353 25087 27387
rect 25087 27353 25096 27387
rect 25044 27344 25096 27353
rect 1768 27319 1820 27328
rect 1768 27285 1777 27319
rect 1777 27285 1811 27319
rect 1811 27285 1820 27319
rect 1768 27276 1820 27285
rect 22836 27319 22888 27328
rect 22836 27285 22845 27319
rect 22845 27285 22879 27319
rect 22879 27285 22888 27319
rect 22836 27276 22888 27285
rect 23480 27276 23532 27328
rect 10214 27174 10266 27226
rect 10278 27174 10330 27226
rect 10342 27174 10394 27226
rect 10406 27174 10458 27226
rect 10470 27174 10522 27226
rect 19478 27174 19530 27226
rect 19542 27174 19594 27226
rect 19606 27174 19658 27226
rect 19670 27174 19722 27226
rect 19734 27174 19786 27226
rect 1676 27072 1728 27124
rect 23480 27115 23532 27124
rect 23480 27081 23489 27115
rect 23489 27081 23523 27115
rect 23523 27081 23532 27115
rect 23480 27072 23532 27081
rect 25136 27115 25188 27124
rect 25136 27081 25145 27115
rect 25145 27081 25179 27115
rect 25179 27081 25188 27115
rect 25136 27072 25188 27081
rect 27528 27072 27580 27124
rect 1400 26979 1452 26988
rect 1400 26945 1409 26979
rect 1409 26945 1443 26979
rect 1443 26945 1452 26979
rect 1400 26936 1452 26945
rect 20904 26868 20956 26920
rect 22376 26979 22428 26988
rect 22376 26945 22410 26979
rect 22410 26945 22428 26979
rect 22376 26936 22428 26945
rect 24032 26979 24084 26988
rect 24032 26945 24066 26979
rect 24066 26945 24084 26979
rect 28080 26979 28132 26988
rect 24032 26936 24084 26945
rect 28080 26945 28089 26979
rect 28089 26945 28123 26979
rect 28123 26945 28132 26979
rect 28080 26936 28132 26945
rect 1584 26775 1636 26784
rect 1584 26741 1593 26775
rect 1593 26741 1627 26775
rect 1627 26741 1636 26775
rect 1584 26732 1636 26741
rect 5582 26630 5634 26682
rect 5646 26630 5698 26682
rect 5710 26630 5762 26682
rect 5774 26630 5826 26682
rect 5838 26630 5890 26682
rect 14846 26630 14898 26682
rect 14910 26630 14962 26682
rect 14974 26630 15026 26682
rect 15038 26630 15090 26682
rect 15102 26630 15154 26682
rect 24110 26630 24162 26682
rect 24174 26630 24226 26682
rect 24238 26630 24290 26682
rect 24302 26630 24354 26682
rect 24366 26630 24418 26682
rect 28356 26571 28408 26580
rect 28356 26537 28365 26571
rect 28365 26537 28399 26571
rect 28399 26537 28408 26571
rect 28356 26528 28408 26537
rect 1400 26367 1452 26376
rect 1400 26333 1409 26367
rect 1409 26333 1443 26367
rect 1443 26333 1452 26367
rect 1400 26324 1452 26333
rect 10214 26086 10266 26138
rect 10278 26086 10330 26138
rect 10342 26086 10394 26138
rect 10406 26086 10458 26138
rect 10470 26086 10522 26138
rect 19478 26086 19530 26138
rect 19542 26086 19594 26138
rect 19606 26086 19658 26138
rect 19670 26086 19722 26138
rect 19734 26086 19786 26138
rect 5582 25542 5634 25594
rect 5646 25542 5698 25594
rect 5710 25542 5762 25594
rect 5774 25542 5826 25594
rect 5838 25542 5890 25594
rect 14846 25542 14898 25594
rect 14910 25542 14962 25594
rect 14974 25542 15026 25594
rect 15038 25542 15090 25594
rect 15102 25542 15154 25594
rect 24110 25542 24162 25594
rect 24174 25542 24226 25594
rect 24238 25542 24290 25594
rect 24302 25542 24354 25594
rect 24366 25542 24418 25594
rect 28356 25279 28408 25288
rect 28356 25245 28365 25279
rect 28365 25245 28399 25279
rect 28399 25245 28408 25279
rect 28356 25236 28408 25245
rect 28172 25143 28224 25152
rect 28172 25109 28181 25143
rect 28181 25109 28215 25143
rect 28215 25109 28224 25143
rect 28172 25100 28224 25109
rect 10214 24998 10266 25050
rect 10278 24998 10330 25050
rect 10342 24998 10394 25050
rect 10406 24998 10458 25050
rect 10470 24998 10522 25050
rect 19478 24998 19530 25050
rect 19542 24998 19594 25050
rect 19606 24998 19658 25050
rect 19670 24998 19722 25050
rect 19734 24998 19786 25050
rect 9036 24828 9088 24880
rect 12164 24828 12216 24880
rect 1400 24803 1452 24812
rect 1400 24769 1409 24803
rect 1409 24769 1443 24803
rect 1443 24769 1452 24803
rect 1400 24760 1452 24769
rect 14740 24760 14792 24812
rect 1676 24556 1728 24608
rect 14648 24556 14700 24608
rect 5582 24454 5634 24506
rect 5646 24454 5698 24506
rect 5710 24454 5762 24506
rect 5774 24454 5826 24506
rect 5838 24454 5890 24506
rect 14846 24454 14898 24506
rect 14910 24454 14962 24506
rect 14974 24454 15026 24506
rect 15038 24454 15090 24506
rect 15102 24454 15154 24506
rect 24110 24454 24162 24506
rect 24174 24454 24226 24506
rect 24238 24454 24290 24506
rect 24302 24454 24354 24506
rect 24366 24454 24418 24506
rect 12900 24148 12952 24200
rect 14648 24191 14700 24200
rect 14648 24157 14682 24191
rect 14682 24157 14700 24191
rect 14648 24148 14700 24157
rect 16304 24148 16356 24200
rect 15568 24012 15620 24064
rect 16396 24012 16448 24064
rect 16948 24012 17000 24064
rect 17224 24055 17276 24064
rect 17224 24021 17233 24055
rect 17233 24021 17267 24055
rect 17267 24021 17276 24055
rect 17224 24012 17276 24021
rect 10214 23910 10266 23962
rect 10278 23910 10330 23962
rect 10342 23910 10394 23962
rect 10406 23910 10458 23962
rect 10470 23910 10522 23962
rect 19478 23910 19530 23962
rect 19542 23910 19594 23962
rect 19606 23910 19658 23962
rect 19670 23910 19722 23962
rect 19734 23910 19786 23962
rect 14740 23808 14792 23860
rect 16304 23851 16356 23860
rect 16304 23817 16313 23851
rect 16313 23817 16347 23851
rect 16347 23817 16356 23851
rect 16304 23808 16356 23817
rect 16396 23808 16448 23860
rect 22836 23808 22888 23860
rect 15292 23783 15344 23792
rect 15292 23749 15301 23783
rect 15301 23749 15335 23783
rect 15335 23749 15344 23783
rect 15292 23740 15344 23749
rect 1400 23511 1452 23520
rect 1400 23477 1409 23511
rect 1409 23477 1443 23511
rect 1443 23477 1452 23511
rect 1400 23468 1452 23477
rect 15568 23672 15620 23724
rect 16120 23715 16172 23724
rect 16120 23681 16129 23715
rect 16129 23681 16163 23715
rect 16163 23681 16172 23715
rect 16120 23672 16172 23681
rect 15476 23647 15528 23656
rect 15476 23613 15485 23647
rect 15485 23613 15519 23647
rect 15519 23613 15528 23647
rect 15476 23604 15528 23613
rect 17132 23740 17184 23792
rect 20904 23783 20956 23792
rect 16948 23715 17000 23724
rect 16948 23681 16982 23715
rect 16982 23681 17000 23715
rect 16948 23672 17000 23681
rect 15660 23468 15712 23520
rect 19248 23536 19300 23588
rect 20904 23749 20913 23783
rect 20913 23749 20947 23783
rect 20947 23749 20956 23783
rect 20904 23740 20956 23749
rect 17040 23468 17092 23520
rect 21180 23468 21232 23520
rect 28356 23511 28408 23520
rect 28356 23477 28365 23511
rect 28365 23477 28399 23511
rect 28399 23477 28408 23511
rect 28356 23468 28408 23477
rect 5582 23366 5634 23418
rect 5646 23366 5698 23418
rect 5710 23366 5762 23418
rect 5774 23366 5826 23418
rect 5838 23366 5890 23418
rect 14846 23366 14898 23418
rect 14910 23366 14962 23418
rect 14974 23366 15026 23418
rect 15038 23366 15090 23418
rect 15102 23366 15154 23418
rect 24110 23366 24162 23418
rect 24174 23366 24226 23418
rect 24238 23366 24290 23418
rect 24302 23366 24354 23418
rect 24366 23366 24418 23418
rect 15292 23307 15344 23316
rect 15292 23273 15301 23307
rect 15301 23273 15335 23307
rect 15335 23273 15344 23307
rect 15292 23264 15344 23273
rect 16120 23264 16172 23316
rect 17224 23264 17276 23316
rect 20536 23264 20588 23316
rect 15476 23196 15528 23248
rect 16488 23196 16540 23248
rect 15660 23128 15712 23180
rect 12624 23060 12676 23112
rect 13452 23103 13504 23112
rect 13452 23069 13461 23103
rect 13461 23069 13495 23103
rect 13495 23069 13504 23103
rect 13452 23060 13504 23069
rect 15752 23103 15804 23112
rect 15752 23069 15761 23103
rect 15761 23069 15795 23103
rect 15795 23069 15804 23103
rect 15752 23060 15804 23069
rect 17224 23060 17276 23112
rect 18420 23103 18472 23112
rect 18420 23069 18429 23103
rect 18429 23069 18463 23103
rect 18463 23069 18472 23103
rect 18420 23060 18472 23069
rect 18880 23103 18932 23112
rect 18880 23069 18889 23103
rect 18889 23069 18923 23103
rect 18923 23069 18932 23103
rect 18880 23060 18932 23069
rect 19984 23060 20036 23112
rect 20260 23103 20312 23112
rect 20260 23069 20269 23103
rect 20269 23069 20303 23103
rect 20303 23069 20312 23103
rect 20260 23060 20312 23069
rect 19248 22992 19300 23044
rect 19340 22992 19392 23044
rect 19892 22992 19944 23044
rect 12992 22967 13044 22976
rect 12992 22933 13001 22967
rect 13001 22933 13035 22967
rect 13035 22933 13044 22967
rect 12992 22924 13044 22933
rect 13268 22967 13320 22976
rect 13268 22933 13277 22967
rect 13277 22933 13311 22967
rect 13311 22933 13320 22967
rect 13268 22924 13320 22933
rect 15568 22924 15620 22976
rect 15844 22924 15896 22976
rect 17040 22924 17092 22976
rect 17132 22924 17184 22976
rect 17960 22967 18012 22976
rect 17960 22933 17969 22967
rect 17969 22933 18003 22967
rect 18003 22933 18012 22967
rect 17960 22924 18012 22933
rect 18236 22967 18288 22976
rect 18236 22933 18245 22967
rect 18245 22933 18279 22967
rect 18279 22933 18288 22967
rect 18236 22924 18288 22933
rect 18696 22967 18748 22976
rect 18696 22933 18705 22967
rect 18705 22933 18739 22967
rect 18739 22933 18748 22967
rect 18696 22924 18748 22933
rect 21456 22924 21508 22976
rect 10214 22822 10266 22874
rect 10278 22822 10330 22874
rect 10342 22822 10394 22874
rect 10406 22822 10458 22874
rect 10470 22822 10522 22874
rect 19478 22822 19530 22874
rect 19542 22822 19594 22874
rect 19606 22822 19658 22874
rect 19670 22822 19722 22874
rect 19734 22822 19786 22874
rect 12624 22763 12676 22772
rect 12624 22729 12633 22763
rect 12633 22729 12667 22763
rect 12667 22729 12676 22763
rect 12624 22720 12676 22729
rect 10876 22584 10928 22636
rect 12532 22652 12584 22704
rect 12992 22652 13044 22704
rect 15292 22652 15344 22704
rect 12900 22627 12952 22636
rect 10508 22423 10560 22432
rect 10508 22389 10517 22423
rect 10517 22389 10551 22423
rect 10551 22389 10560 22423
rect 10508 22380 10560 22389
rect 12900 22593 12909 22627
rect 12909 22593 12943 22627
rect 12943 22593 12952 22627
rect 12900 22584 12952 22593
rect 15844 22720 15896 22772
rect 17224 22720 17276 22772
rect 17132 22652 17184 22704
rect 15844 22627 15896 22636
rect 15844 22593 15853 22627
rect 15853 22593 15887 22627
rect 15887 22593 15896 22627
rect 15844 22584 15896 22593
rect 15936 22627 15988 22636
rect 15936 22593 15945 22627
rect 15945 22593 15979 22627
rect 15979 22593 15988 22627
rect 15936 22584 15988 22593
rect 17960 22584 18012 22636
rect 18696 22652 18748 22704
rect 20904 22652 20956 22704
rect 14188 22516 14240 22568
rect 19340 22584 19392 22636
rect 20628 22584 20680 22636
rect 21364 22584 21416 22636
rect 13912 22448 13964 22500
rect 15844 22448 15896 22500
rect 16672 22423 16724 22432
rect 16672 22389 16681 22423
rect 16681 22389 16715 22423
rect 16715 22389 16724 22423
rect 16672 22380 16724 22389
rect 19064 22380 19116 22432
rect 19708 22423 19760 22432
rect 19708 22389 19717 22423
rect 19717 22389 19751 22423
rect 19751 22389 19760 22423
rect 19708 22380 19760 22389
rect 5582 22278 5634 22330
rect 5646 22278 5698 22330
rect 5710 22278 5762 22330
rect 5774 22278 5826 22330
rect 5838 22278 5890 22330
rect 14846 22278 14898 22330
rect 14910 22278 14962 22330
rect 14974 22278 15026 22330
rect 15038 22278 15090 22330
rect 15102 22278 15154 22330
rect 24110 22278 24162 22330
rect 24174 22278 24226 22330
rect 24238 22278 24290 22330
rect 24302 22278 24354 22330
rect 24366 22278 24418 22330
rect 15752 22176 15804 22228
rect 16672 22176 16724 22228
rect 17592 22176 17644 22228
rect 18880 22219 18932 22228
rect 18880 22185 18889 22219
rect 18889 22185 18923 22219
rect 18923 22185 18932 22219
rect 18880 22176 18932 22185
rect 20260 22219 20312 22228
rect 20260 22185 20269 22219
rect 20269 22185 20303 22219
rect 20303 22185 20312 22219
rect 20260 22176 20312 22185
rect 21364 22176 21416 22228
rect 16488 22108 16540 22160
rect 16304 22040 16356 22092
rect 7564 21972 7616 22024
rect 9680 21972 9732 22024
rect 10508 21972 10560 22024
rect 12440 21972 12492 22024
rect 12900 21972 12952 22024
rect 17132 21972 17184 22024
rect 17224 21972 17276 22024
rect 18788 22108 18840 22160
rect 19064 22108 19116 22160
rect 17592 21972 17644 22024
rect 18972 22040 19024 22092
rect 19892 22083 19944 22092
rect 19892 22049 19901 22083
rect 19901 22049 19935 22083
rect 19935 22049 19944 22083
rect 19892 22040 19944 22049
rect 18604 22015 18656 22024
rect 10140 21947 10192 21956
rect 10140 21913 10149 21947
rect 10149 21913 10183 21947
rect 10183 21913 10192 21947
rect 10140 21904 10192 21913
rect 11612 21904 11664 21956
rect 13268 21904 13320 21956
rect 16488 21904 16540 21956
rect 7932 21836 7984 21888
rect 9404 21879 9456 21888
rect 9404 21845 9413 21879
rect 9413 21845 9447 21879
rect 9447 21845 9456 21879
rect 9404 21836 9456 21845
rect 12716 21836 12768 21888
rect 13912 21836 13964 21888
rect 14004 21836 14056 21888
rect 16580 21879 16632 21888
rect 16580 21845 16589 21879
rect 16589 21845 16623 21879
rect 16623 21845 16632 21879
rect 16580 21836 16632 21845
rect 16672 21879 16724 21888
rect 16672 21845 16681 21879
rect 16681 21845 16715 21879
rect 16715 21845 16724 21879
rect 16672 21836 16724 21845
rect 17040 21836 17092 21888
rect 18604 21981 18613 22015
rect 18613 21981 18647 22015
rect 18647 21981 18656 22015
rect 18604 21972 18656 21981
rect 18696 22015 18748 22024
rect 18696 21981 18705 22015
rect 18705 21981 18739 22015
rect 18739 21981 18748 22015
rect 18696 21972 18748 21981
rect 20536 21972 20588 22024
rect 18788 21904 18840 21956
rect 19708 21947 19760 21956
rect 19708 21913 19717 21947
rect 19717 21913 19751 21947
rect 19751 21913 19760 21947
rect 19708 21904 19760 21913
rect 19892 21904 19944 21956
rect 21456 22015 21508 22024
rect 21456 21981 21465 22015
rect 21465 21981 21499 22015
rect 21499 21981 21508 22015
rect 21456 21972 21508 21981
rect 17960 21879 18012 21888
rect 17960 21845 17969 21879
rect 17969 21845 18003 21879
rect 18003 21845 18012 21879
rect 17960 21836 18012 21845
rect 18696 21836 18748 21888
rect 19340 21836 19392 21888
rect 10214 21734 10266 21786
rect 10278 21734 10330 21786
rect 10342 21734 10394 21786
rect 10406 21734 10458 21786
rect 10470 21734 10522 21786
rect 19478 21734 19530 21786
rect 19542 21734 19594 21786
rect 19606 21734 19658 21786
rect 19670 21734 19722 21786
rect 19734 21734 19786 21786
rect 9772 21632 9824 21684
rect 13452 21632 13504 21684
rect 13912 21632 13964 21684
rect 16488 21632 16540 21684
rect 18420 21632 18472 21684
rect 20536 21632 20588 21684
rect 25044 21632 25096 21684
rect 6828 21496 6880 21548
rect 7932 21539 7984 21548
rect 7932 21505 7966 21539
rect 7966 21505 7984 21539
rect 7932 21496 7984 21505
rect 9404 21564 9456 21616
rect 12624 21564 12676 21616
rect 11152 21496 11204 21548
rect 15292 21564 15344 21616
rect 9128 21428 9180 21480
rect 12348 21428 12400 21480
rect 12532 21471 12584 21480
rect 12532 21437 12541 21471
rect 12541 21437 12575 21471
rect 12575 21437 12584 21471
rect 12532 21428 12584 21437
rect 1400 21335 1452 21344
rect 1400 21301 1409 21335
rect 1409 21301 1443 21335
rect 1443 21301 1452 21335
rect 1400 21292 1452 21301
rect 7656 21292 7708 21344
rect 9036 21335 9088 21344
rect 9036 21301 9045 21335
rect 9045 21301 9079 21335
rect 9079 21301 9088 21335
rect 9036 21292 9088 21301
rect 11336 21292 11388 21344
rect 11520 21335 11572 21344
rect 11520 21301 11529 21335
rect 11529 21301 11563 21335
rect 11563 21301 11572 21335
rect 11520 21292 11572 21301
rect 13452 21292 13504 21344
rect 14004 21496 14056 21548
rect 15844 21496 15896 21548
rect 14188 21471 14240 21480
rect 14188 21437 14197 21471
rect 14197 21437 14231 21471
rect 14231 21437 14240 21471
rect 14188 21428 14240 21437
rect 15752 21471 15804 21480
rect 15752 21437 15761 21471
rect 15761 21437 15795 21471
rect 15795 21437 15804 21471
rect 15752 21428 15804 21437
rect 17132 21496 17184 21548
rect 18236 21564 18288 21616
rect 18604 21564 18656 21616
rect 18880 21496 18932 21548
rect 19616 21496 19668 21548
rect 19984 21539 20036 21548
rect 19984 21505 19993 21539
rect 19993 21505 20027 21539
rect 20027 21505 20036 21539
rect 19984 21496 20036 21505
rect 20168 21539 20220 21548
rect 20168 21505 20177 21539
rect 20177 21505 20211 21539
rect 20211 21505 20220 21539
rect 20168 21496 20220 21505
rect 20260 21496 20312 21548
rect 19984 21360 20036 21412
rect 15568 21292 15620 21344
rect 16580 21292 16632 21344
rect 17224 21335 17276 21344
rect 17224 21301 17233 21335
rect 17233 21301 17267 21335
rect 17267 21301 17276 21335
rect 17224 21292 17276 21301
rect 18420 21292 18472 21344
rect 20904 21292 20956 21344
rect 21272 21292 21324 21344
rect 5582 21190 5634 21242
rect 5646 21190 5698 21242
rect 5710 21190 5762 21242
rect 5774 21190 5826 21242
rect 5838 21190 5890 21242
rect 14846 21190 14898 21242
rect 14910 21190 14962 21242
rect 14974 21190 15026 21242
rect 15038 21190 15090 21242
rect 15102 21190 15154 21242
rect 24110 21190 24162 21242
rect 24174 21190 24226 21242
rect 24238 21190 24290 21242
rect 24302 21190 24354 21242
rect 24366 21190 24418 21242
rect 7564 21131 7616 21140
rect 7564 21097 7573 21131
rect 7573 21097 7607 21131
rect 7607 21097 7616 21131
rect 7564 21088 7616 21097
rect 11612 21131 11664 21140
rect 3148 21020 3200 21072
rect 7656 21020 7708 21072
rect 11612 21097 11621 21131
rect 11621 21097 11655 21131
rect 11655 21097 11664 21131
rect 11612 21088 11664 21097
rect 15752 21088 15804 21140
rect 18880 21131 18932 21140
rect 9404 21020 9456 21072
rect 8116 20952 8168 21004
rect 8208 20884 8260 20936
rect 9772 20927 9824 20936
rect 9772 20893 9781 20927
rect 9781 20893 9815 20927
rect 9815 20893 9824 20927
rect 9772 20884 9824 20893
rect 10876 20927 10928 20936
rect 10876 20893 10885 20927
rect 10885 20893 10919 20927
rect 10919 20893 10928 20927
rect 10876 20884 10928 20893
rect 11520 20952 11572 21004
rect 16764 21020 16816 21072
rect 16304 20995 16356 21004
rect 16304 20961 16313 20995
rect 16313 20961 16347 20995
rect 16347 20961 16356 20995
rect 16304 20952 16356 20961
rect 12440 20884 12492 20936
rect 13544 20884 13596 20936
rect 15292 20927 15344 20936
rect 15292 20893 15301 20927
rect 15301 20893 15335 20927
rect 15335 20893 15344 20927
rect 15292 20884 15344 20893
rect 18880 21097 18889 21131
rect 18889 21097 18923 21131
rect 18923 21097 18932 21131
rect 18880 21088 18932 21097
rect 20260 21088 20312 21140
rect 28080 21088 28132 21140
rect 18420 20995 18472 21004
rect 9036 20816 9088 20868
rect 11244 20816 11296 20868
rect 11336 20816 11388 20868
rect 18420 20961 18429 20995
rect 18429 20961 18463 20995
rect 18463 20961 18472 20995
rect 18420 20952 18472 20961
rect 19340 20995 19392 21004
rect 19340 20961 19349 20995
rect 19349 20961 19383 20995
rect 19383 20961 19392 20995
rect 19340 20952 19392 20961
rect 19616 20952 19668 21004
rect 21272 20884 21324 20936
rect 23204 20884 23256 20936
rect 19892 20816 19944 20868
rect 20536 20816 20588 20868
rect 22468 20816 22520 20868
rect 9496 20748 9548 20800
rect 12808 20748 12860 20800
rect 13452 20748 13504 20800
rect 16120 20748 16172 20800
rect 19248 20748 19300 20800
rect 20260 20748 20312 20800
rect 20444 20791 20496 20800
rect 20444 20757 20453 20791
rect 20453 20757 20487 20791
rect 20487 20757 20496 20791
rect 20444 20748 20496 20757
rect 10214 20646 10266 20698
rect 10278 20646 10330 20698
rect 10342 20646 10394 20698
rect 10406 20646 10458 20698
rect 10470 20646 10522 20698
rect 19478 20646 19530 20698
rect 19542 20646 19594 20698
rect 19606 20646 19658 20698
rect 19670 20646 19722 20698
rect 19734 20646 19786 20698
rect 9680 20587 9732 20596
rect 9680 20553 9689 20587
rect 9689 20553 9723 20587
rect 9723 20553 9732 20587
rect 9680 20544 9732 20553
rect 11152 20587 11204 20596
rect 11152 20553 11161 20587
rect 11161 20553 11195 20587
rect 11195 20553 11204 20587
rect 11152 20544 11204 20553
rect 11244 20544 11296 20596
rect 15476 20544 15528 20596
rect 10140 20476 10192 20528
rect 7104 20451 7156 20460
rect 7104 20417 7138 20451
rect 7138 20417 7156 20451
rect 9496 20451 9548 20460
rect 7104 20408 7156 20417
rect 9496 20417 9505 20451
rect 9505 20417 9539 20451
rect 9539 20417 9548 20451
rect 9496 20408 9548 20417
rect 10048 20408 10100 20460
rect 10876 20451 10928 20460
rect 10876 20417 10885 20451
rect 10885 20417 10919 20451
rect 10919 20417 10928 20451
rect 10876 20408 10928 20417
rect 6828 20383 6880 20392
rect 6828 20349 6837 20383
rect 6837 20349 6871 20383
rect 6871 20349 6880 20383
rect 6828 20340 6880 20349
rect 9404 20340 9456 20392
rect 12808 20408 12860 20460
rect 13636 20408 13688 20460
rect 14280 20451 14332 20460
rect 14280 20417 14289 20451
rect 14289 20417 14323 20451
rect 14323 20417 14332 20451
rect 14280 20408 14332 20417
rect 15568 20408 15620 20460
rect 12348 20383 12400 20392
rect 12348 20349 12357 20383
rect 12357 20349 12391 20383
rect 12391 20349 12400 20383
rect 12348 20340 12400 20349
rect 16304 20476 16356 20528
rect 17132 20476 17184 20528
rect 18328 20544 18380 20596
rect 19340 20544 19392 20596
rect 20168 20544 20220 20596
rect 16764 20408 16816 20460
rect 18788 20451 18840 20460
rect 18788 20417 18797 20451
rect 18797 20417 18831 20451
rect 18831 20417 18840 20451
rect 20444 20476 20496 20528
rect 18788 20408 18840 20417
rect 19156 20451 19208 20460
rect 19156 20417 19165 20451
rect 19165 20417 19199 20451
rect 19199 20417 19208 20451
rect 19156 20408 19208 20417
rect 19984 20408 20036 20460
rect 20168 20408 20220 20460
rect 20904 20451 20956 20460
rect 20904 20417 20913 20451
rect 20913 20417 20947 20451
rect 20947 20417 20956 20451
rect 20904 20408 20956 20417
rect 20536 20383 20588 20392
rect 13544 20272 13596 20324
rect 20536 20349 20545 20383
rect 20545 20349 20579 20383
rect 20579 20349 20588 20383
rect 20536 20340 20588 20349
rect 23204 20383 23256 20392
rect 23204 20349 23213 20383
rect 23213 20349 23247 20383
rect 23247 20349 23256 20383
rect 23204 20340 23256 20349
rect 8208 20247 8260 20256
rect 8208 20213 8217 20247
rect 8217 20213 8251 20247
rect 8251 20213 8260 20247
rect 8208 20204 8260 20213
rect 9128 20204 9180 20256
rect 11704 20204 11756 20256
rect 13912 20247 13964 20256
rect 13912 20213 13921 20247
rect 13921 20213 13955 20247
rect 13955 20213 13964 20247
rect 13912 20204 13964 20213
rect 14556 20247 14608 20256
rect 14556 20213 14565 20247
rect 14565 20213 14599 20247
rect 14599 20213 14608 20247
rect 14556 20204 14608 20213
rect 16120 20204 16172 20256
rect 18420 20204 18472 20256
rect 5582 20102 5634 20154
rect 5646 20102 5698 20154
rect 5710 20102 5762 20154
rect 5774 20102 5826 20154
rect 5838 20102 5890 20154
rect 14846 20102 14898 20154
rect 14910 20102 14962 20154
rect 14974 20102 15026 20154
rect 15038 20102 15090 20154
rect 15102 20102 15154 20154
rect 24110 20102 24162 20154
rect 24174 20102 24226 20154
rect 24238 20102 24290 20154
rect 24302 20102 24354 20154
rect 24366 20102 24418 20154
rect 7104 20000 7156 20052
rect 12348 20000 12400 20052
rect 15476 20043 15528 20052
rect 1400 19839 1452 19848
rect 1400 19805 1409 19839
rect 1409 19805 1443 19839
rect 1443 19805 1452 19839
rect 1400 19796 1452 19805
rect 8116 19864 8168 19916
rect 13544 19864 13596 19916
rect 15476 20009 15485 20043
rect 15485 20009 15519 20043
rect 15519 20009 15528 20043
rect 15476 20000 15528 20009
rect 16212 20000 16264 20052
rect 19156 20000 19208 20052
rect 19248 20000 19300 20052
rect 22744 20000 22796 20052
rect 20076 19932 20128 19984
rect 8300 19796 8352 19848
rect 9036 19839 9088 19848
rect 9036 19805 9045 19839
rect 9045 19805 9079 19839
rect 9079 19805 9088 19839
rect 9036 19796 9088 19805
rect 9128 19796 9180 19848
rect 13084 19796 13136 19848
rect 7748 19728 7800 19780
rect 9312 19771 9364 19780
rect 9312 19737 9346 19771
rect 9346 19737 9364 19771
rect 9312 19728 9364 19737
rect 11520 19728 11572 19780
rect 13912 19796 13964 19848
rect 16120 19839 16172 19848
rect 15292 19728 15344 19780
rect 16120 19805 16129 19839
rect 16129 19805 16163 19839
rect 16163 19805 16172 19839
rect 16120 19796 16172 19805
rect 16580 19796 16632 19848
rect 17684 19796 17736 19848
rect 17960 19839 18012 19848
rect 17960 19805 17969 19839
rect 17969 19805 18003 19839
rect 18003 19805 18012 19839
rect 17960 19796 18012 19805
rect 19892 19864 19944 19916
rect 20260 19864 20312 19916
rect 22100 19864 22152 19916
rect 18328 19839 18380 19848
rect 18328 19805 18337 19839
rect 18337 19805 18371 19839
rect 18371 19805 18380 19839
rect 18328 19796 18380 19805
rect 18420 19839 18472 19848
rect 18420 19805 18434 19839
rect 18434 19805 18468 19839
rect 18468 19805 18472 19839
rect 18420 19796 18472 19805
rect 20628 19796 20680 19848
rect 24216 19796 24268 19848
rect 8208 19703 8260 19712
rect 8208 19669 8217 19703
rect 8217 19669 8251 19703
rect 8251 19669 8260 19703
rect 8208 19660 8260 19669
rect 9680 19660 9732 19712
rect 12256 19660 12308 19712
rect 14280 19660 14332 19712
rect 15752 19703 15804 19712
rect 15752 19669 15761 19703
rect 15761 19669 15795 19703
rect 15795 19669 15804 19703
rect 15752 19660 15804 19669
rect 16028 19728 16080 19780
rect 18236 19771 18288 19780
rect 17408 19660 17460 19712
rect 18236 19737 18245 19771
rect 18245 19737 18279 19771
rect 18279 19737 18288 19771
rect 18236 19728 18288 19737
rect 20260 19728 20312 19780
rect 20168 19660 20220 19712
rect 20536 19703 20588 19712
rect 20536 19669 20545 19703
rect 20545 19669 20579 19703
rect 20579 19669 20588 19703
rect 20536 19660 20588 19669
rect 21088 19703 21140 19712
rect 21088 19669 21097 19703
rect 21097 19669 21131 19703
rect 21131 19669 21140 19703
rect 21732 19728 21784 19780
rect 22652 19771 22704 19780
rect 22652 19737 22686 19771
rect 22686 19737 22704 19771
rect 22652 19728 22704 19737
rect 21088 19660 21140 19669
rect 23020 19660 23072 19712
rect 10214 19558 10266 19610
rect 10278 19558 10330 19610
rect 10342 19558 10394 19610
rect 10406 19558 10458 19610
rect 10470 19558 10522 19610
rect 19478 19558 19530 19610
rect 19542 19558 19594 19610
rect 19606 19558 19658 19610
rect 19670 19558 19722 19610
rect 19734 19558 19786 19610
rect 1400 19499 1452 19508
rect 1400 19465 1409 19499
rect 1409 19465 1443 19499
rect 1443 19465 1452 19499
rect 1400 19456 1452 19465
rect 6920 19456 6972 19508
rect 9312 19499 9364 19508
rect 9312 19465 9321 19499
rect 9321 19465 9355 19499
rect 9355 19465 9364 19499
rect 9312 19456 9364 19465
rect 10048 19456 10100 19508
rect 11520 19499 11572 19508
rect 11520 19465 11529 19499
rect 11529 19465 11563 19499
rect 11563 19465 11572 19499
rect 11520 19456 11572 19465
rect 13636 19499 13688 19508
rect 13636 19465 13645 19499
rect 13645 19465 13679 19499
rect 13679 19465 13688 19499
rect 13636 19456 13688 19465
rect 15476 19499 15528 19508
rect 15476 19465 15485 19499
rect 15485 19465 15519 19499
rect 15519 19465 15528 19499
rect 15476 19456 15528 19465
rect 16212 19499 16264 19508
rect 16212 19465 16221 19499
rect 16221 19465 16255 19499
rect 16255 19465 16264 19499
rect 16212 19456 16264 19465
rect 8208 19388 8260 19440
rect 7012 19363 7064 19372
rect 7012 19329 7021 19363
rect 7021 19329 7055 19363
rect 7055 19329 7064 19363
rect 7012 19320 7064 19329
rect 8852 19363 8904 19372
rect 8852 19329 8861 19363
rect 8861 19329 8895 19363
rect 8895 19329 8904 19363
rect 8852 19320 8904 19329
rect 12256 19388 12308 19440
rect 17040 19499 17092 19508
rect 17040 19465 17049 19499
rect 17049 19465 17083 19499
rect 17083 19465 17092 19499
rect 17040 19456 17092 19465
rect 18788 19456 18840 19508
rect 20444 19456 20496 19508
rect 11704 19363 11756 19372
rect 11704 19329 11713 19363
rect 11713 19329 11747 19363
rect 11747 19329 11756 19363
rect 11704 19320 11756 19329
rect 12532 19320 12584 19372
rect 14556 19320 14608 19372
rect 16028 19363 16080 19372
rect 8300 19252 8352 19304
rect 9404 19252 9456 19304
rect 10968 19295 11020 19304
rect 10968 19261 10977 19295
rect 10977 19261 11011 19295
rect 11011 19261 11020 19295
rect 10968 19252 11020 19261
rect 11244 19252 11296 19304
rect 13084 19252 13136 19304
rect 14648 19252 14700 19304
rect 16028 19329 16037 19363
rect 16037 19329 16071 19363
rect 16071 19329 16080 19363
rect 16028 19320 16080 19329
rect 16580 19320 16632 19372
rect 19340 19388 19392 19440
rect 19616 19388 19668 19440
rect 22652 19456 22704 19508
rect 24216 19431 24268 19440
rect 24216 19397 24225 19431
rect 24225 19397 24259 19431
rect 24259 19397 24268 19431
rect 24216 19388 24268 19397
rect 17776 19363 17828 19372
rect 17776 19329 17810 19363
rect 17810 19329 17828 19363
rect 17776 19320 17828 19329
rect 20076 19320 20128 19372
rect 20628 19363 20680 19372
rect 20628 19329 20637 19363
rect 20637 19329 20671 19363
rect 20671 19329 20680 19363
rect 20628 19320 20680 19329
rect 20812 19320 20864 19372
rect 21732 19320 21784 19372
rect 20904 19252 20956 19304
rect 22304 19363 22356 19372
rect 22304 19329 22313 19363
rect 22313 19329 22347 19363
rect 22347 19329 22356 19363
rect 23020 19363 23072 19372
rect 22304 19320 22356 19329
rect 23020 19329 23029 19363
rect 23029 19329 23063 19363
rect 23063 19329 23072 19363
rect 23020 19320 23072 19329
rect 23296 19320 23348 19372
rect 23664 19363 23716 19372
rect 23664 19329 23673 19363
rect 23673 19329 23707 19363
rect 23707 19329 23716 19363
rect 23664 19320 23716 19329
rect 22652 19252 22704 19304
rect 23572 19252 23624 19304
rect 24676 19295 24728 19304
rect 24676 19261 24685 19295
rect 24685 19261 24719 19295
rect 24719 19261 24728 19295
rect 24676 19252 24728 19261
rect 1584 19116 1636 19168
rect 11336 19184 11388 19236
rect 14096 19184 14148 19236
rect 14740 19116 14792 19168
rect 15292 19116 15344 19168
rect 15936 19116 15988 19168
rect 16764 19116 16816 19168
rect 19616 19116 19668 19168
rect 23204 19184 23256 19236
rect 20720 19116 20772 19168
rect 21456 19159 21508 19168
rect 21456 19125 21465 19159
rect 21465 19125 21499 19159
rect 21499 19125 21508 19159
rect 21456 19116 21508 19125
rect 23848 19159 23900 19168
rect 23848 19125 23857 19159
rect 23857 19125 23891 19159
rect 23891 19125 23900 19159
rect 23848 19116 23900 19125
rect 23940 19116 23992 19168
rect 5582 19014 5634 19066
rect 5646 19014 5698 19066
rect 5710 19014 5762 19066
rect 5774 19014 5826 19066
rect 5838 19014 5890 19066
rect 14846 19014 14898 19066
rect 14910 19014 14962 19066
rect 14974 19014 15026 19066
rect 15038 19014 15090 19066
rect 15102 19014 15154 19066
rect 24110 19014 24162 19066
rect 24174 19014 24226 19066
rect 24238 19014 24290 19066
rect 24302 19014 24354 19066
rect 24366 19014 24418 19066
rect 8852 18912 8904 18964
rect 10876 18912 10928 18964
rect 1400 18751 1452 18760
rect 1400 18717 1409 18751
rect 1409 18717 1443 18751
rect 1443 18717 1452 18751
rect 1400 18708 1452 18717
rect 6644 18751 6696 18760
rect 6644 18717 6653 18751
rect 6653 18717 6687 18751
rect 6687 18717 6696 18751
rect 6644 18708 6696 18717
rect 6920 18751 6972 18760
rect 6920 18717 6954 18751
rect 6954 18717 6972 18751
rect 6920 18708 6972 18717
rect 7288 18708 7340 18760
rect 8116 18776 8168 18828
rect 10968 18819 11020 18828
rect 10968 18785 10977 18819
rect 10977 18785 11011 18819
rect 11011 18785 11020 18819
rect 10968 18776 11020 18785
rect 9680 18708 9732 18760
rect 7840 18572 7892 18624
rect 9588 18640 9640 18692
rect 12716 18912 12768 18964
rect 14372 18912 14424 18964
rect 16764 18912 16816 18964
rect 17776 18912 17828 18964
rect 19340 18912 19392 18964
rect 20628 18912 20680 18964
rect 20720 18912 20772 18964
rect 13820 18844 13872 18896
rect 12256 18683 12308 18692
rect 12256 18649 12265 18683
rect 12265 18649 12299 18683
rect 12299 18649 12308 18683
rect 12256 18640 12308 18649
rect 10692 18572 10744 18624
rect 11428 18572 11480 18624
rect 11612 18615 11664 18624
rect 11612 18581 11621 18615
rect 11621 18581 11655 18615
rect 11655 18581 11664 18615
rect 11612 18572 11664 18581
rect 12440 18615 12492 18624
rect 12440 18581 12465 18615
rect 12465 18581 12492 18615
rect 12808 18640 12860 18692
rect 14188 18708 14240 18760
rect 14372 18751 14424 18760
rect 14372 18717 14381 18751
rect 14381 18717 14415 18751
rect 14415 18717 14424 18751
rect 14372 18708 14424 18717
rect 14556 18844 14608 18896
rect 14740 18844 14792 18896
rect 15108 18819 15160 18828
rect 14648 18708 14700 18760
rect 15108 18785 15117 18819
rect 15117 18785 15151 18819
rect 15151 18785 15160 18819
rect 15108 18776 15160 18785
rect 17316 18776 17368 18828
rect 14832 18708 14884 18760
rect 15292 18751 15344 18760
rect 15292 18717 15301 18751
rect 15301 18717 15335 18751
rect 15335 18717 15344 18751
rect 15292 18708 15344 18717
rect 12440 18572 12492 18581
rect 14004 18572 14056 18624
rect 16028 18708 16080 18760
rect 16580 18708 16632 18760
rect 16948 18708 17000 18760
rect 17408 18751 17460 18760
rect 16672 18640 16724 18692
rect 17408 18717 17417 18751
rect 17417 18717 17451 18751
rect 17451 18717 17460 18751
rect 17408 18708 17460 18717
rect 17776 18776 17828 18828
rect 17684 18708 17736 18760
rect 17960 18708 18012 18760
rect 18144 18751 18196 18760
rect 18144 18717 18153 18751
rect 18153 18717 18187 18751
rect 18187 18717 18196 18751
rect 18144 18708 18196 18717
rect 20260 18708 20312 18760
rect 20720 18751 20772 18760
rect 15660 18572 15712 18624
rect 16212 18572 16264 18624
rect 19248 18640 19300 18692
rect 19616 18683 19668 18692
rect 19616 18649 19625 18683
rect 19625 18649 19659 18683
rect 19659 18649 19668 18683
rect 19616 18640 19668 18649
rect 20168 18640 20220 18692
rect 18052 18572 18104 18624
rect 18328 18615 18380 18624
rect 18328 18581 18337 18615
rect 18337 18581 18371 18615
rect 18371 18581 18380 18615
rect 18328 18572 18380 18581
rect 20076 18615 20128 18624
rect 20076 18581 20085 18615
rect 20085 18581 20119 18615
rect 20119 18581 20128 18615
rect 20076 18572 20128 18581
rect 20720 18717 20729 18751
rect 20729 18717 20763 18751
rect 20763 18717 20772 18751
rect 20720 18708 20772 18717
rect 21180 18708 21232 18760
rect 21456 18751 21508 18760
rect 20628 18640 20680 18692
rect 20536 18572 20588 18624
rect 21456 18717 21465 18751
rect 21465 18717 21499 18751
rect 21499 18717 21508 18751
rect 21456 18708 21508 18717
rect 22376 18912 22428 18964
rect 23664 18912 23716 18964
rect 21824 18844 21876 18896
rect 22284 18708 22336 18760
rect 22928 18708 22980 18760
rect 23848 18776 23900 18828
rect 23480 18751 23532 18760
rect 23480 18717 23510 18751
rect 23510 18717 23532 18751
rect 23480 18708 23532 18717
rect 23572 18751 23624 18760
rect 23572 18717 23601 18751
rect 23601 18717 23624 18751
rect 23572 18708 23624 18717
rect 23940 18708 23992 18760
rect 21732 18640 21784 18692
rect 21824 18572 21876 18624
rect 22008 18572 22060 18624
rect 22652 18572 22704 18624
rect 23480 18572 23532 18624
rect 10214 18470 10266 18522
rect 10278 18470 10330 18522
rect 10342 18470 10394 18522
rect 10406 18470 10458 18522
rect 10470 18470 10522 18522
rect 19478 18470 19530 18522
rect 19542 18470 19594 18522
rect 19606 18470 19658 18522
rect 19670 18470 19722 18522
rect 19734 18470 19786 18522
rect 7012 18368 7064 18420
rect 7840 18411 7892 18420
rect 6000 18207 6052 18216
rect 6000 18173 6009 18207
rect 6009 18173 6043 18207
rect 6043 18173 6052 18207
rect 6000 18164 6052 18173
rect 6736 18207 6788 18216
rect 6736 18173 6745 18207
rect 6745 18173 6779 18207
rect 6779 18173 6788 18207
rect 6736 18164 6788 18173
rect 7840 18377 7849 18411
rect 7849 18377 7883 18411
rect 7883 18377 7892 18411
rect 7840 18368 7892 18377
rect 7288 18164 7340 18216
rect 7380 18164 7432 18216
rect 8116 18207 8168 18216
rect 8116 18173 8125 18207
rect 8125 18173 8159 18207
rect 8159 18173 8168 18207
rect 8116 18164 8168 18173
rect 6644 18096 6696 18148
rect 9036 18368 9088 18420
rect 9588 18411 9640 18420
rect 9588 18377 9597 18411
rect 9597 18377 9631 18411
rect 9631 18377 9640 18411
rect 9588 18368 9640 18377
rect 9680 18368 9732 18420
rect 10968 18368 11020 18420
rect 11428 18368 11480 18420
rect 13820 18411 13872 18420
rect 9864 18300 9916 18352
rect 10324 18232 10376 18284
rect 9680 18207 9732 18216
rect 9680 18173 9689 18207
rect 9689 18173 9723 18207
rect 9723 18173 9732 18207
rect 9680 18164 9732 18173
rect 9772 18164 9824 18216
rect 4620 18071 4672 18080
rect 4620 18037 4629 18071
rect 4629 18037 4663 18071
rect 4663 18037 4672 18071
rect 4620 18028 4672 18037
rect 6736 18028 6788 18080
rect 9128 18071 9180 18080
rect 9128 18037 9137 18071
rect 9137 18037 9171 18071
rect 9171 18037 9180 18071
rect 9128 18028 9180 18037
rect 13084 18300 13136 18352
rect 13820 18377 13829 18411
rect 13829 18377 13863 18411
rect 13863 18377 13872 18411
rect 13820 18368 13872 18377
rect 14648 18368 14700 18420
rect 13544 18300 13596 18352
rect 10692 18232 10744 18284
rect 11152 18232 11204 18284
rect 14004 18275 14056 18284
rect 14004 18241 14013 18275
rect 14013 18241 14047 18275
rect 14047 18241 14056 18275
rect 14004 18232 14056 18241
rect 14096 18275 14148 18284
rect 14096 18241 14105 18275
rect 14105 18241 14139 18275
rect 14139 18241 14148 18275
rect 14372 18275 14424 18284
rect 14096 18232 14148 18241
rect 14372 18241 14381 18275
rect 14381 18241 14415 18275
rect 14415 18241 14424 18275
rect 14372 18232 14424 18241
rect 15752 18300 15804 18352
rect 17040 18300 17092 18352
rect 17316 18300 17368 18352
rect 11520 18207 11572 18216
rect 11520 18173 11529 18207
rect 11529 18173 11563 18207
rect 11563 18173 11572 18207
rect 11520 18164 11572 18173
rect 15292 18232 15344 18284
rect 16028 18275 16080 18284
rect 16028 18241 16037 18275
rect 16037 18241 16071 18275
rect 16071 18241 16080 18275
rect 16028 18232 16080 18241
rect 16948 18275 17000 18284
rect 16948 18241 16957 18275
rect 16957 18241 16991 18275
rect 16991 18241 17000 18275
rect 16948 18232 17000 18241
rect 19340 18300 19392 18352
rect 19892 18368 19944 18420
rect 20168 18368 20220 18420
rect 20444 18343 20496 18352
rect 20444 18309 20453 18343
rect 20453 18309 20487 18343
rect 20487 18309 20496 18343
rect 20444 18300 20496 18309
rect 18328 18232 18380 18284
rect 19248 18232 19300 18284
rect 20720 18300 20772 18352
rect 20904 18300 20956 18352
rect 22100 18368 22152 18420
rect 22468 18411 22520 18420
rect 22468 18377 22477 18411
rect 22477 18377 22511 18411
rect 22511 18377 22520 18411
rect 22468 18368 22520 18377
rect 21916 18300 21968 18352
rect 20812 18232 20864 18284
rect 21088 18275 21140 18284
rect 21088 18241 21097 18275
rect 21097 18241 21131 18275
rect 21131 18241 21140 18275
rect 21088 18232 21140 18241
rect 21824 18275 21876 18284
rect 21824 18241 21833 18275
rect 21833 18241 21867 18275
rect 21867 18241 21876 18275
rect 21824 18232 21876 18241
rect 22008 18275 22060 18284
rect 22008 18241 22017 18275
rect 22017 18241 22051 18275
rect 22051 18241 22060 18275
rect 22008 18232 22060 18241
rect 22744 18300 22796 18352
rect 22284 18232 22336 18284
rect 23020 18275 23072 18284
rect 23020 18241 23024 18275
rect 23024 18241 23058 18275
rect 23058 18241 23072 18275
rect 15108 18207 15160 18216
rect 15108 18173 15117 18207
rect 15117 18173 15151 18207
rect 15151 18173 15160 18207
rect 15108 18164 15160 18173
rect 15476 18164 15528 18216
rect 16396 18164 16448 18216
rect 16672 18207 16724 18216
rect 16672 18173 16681 18207
rect 16681 18173 16715 18207
rect 16715 18173 16724 18207
rect 16672 18164 16724 18173
rect 10968 18028 11020 18080
rect 13360 18071 13412 18080
rect 13360 18037 13369 18071
rect 13369 18037 13403 18071
rect 13403 18037 13412 18071
rect 13360 18028 13412 18037
rect 14464 18028 14516 18080
rect 18052 18028 18104 18080
rect 20536 18096 20588 18148
rect 20628 18096 20680 18148
rect 22652 18096 22704 18148
rect 20444 18028 20496 18080
rect 20720 18028 20772 18080
rect 23020 18232 23072 18241
rect 23848 18232 23900 18284
rect 23480 18164 23532 18216
rect 22928 18028 22980 18080
rect 23112 18028 23164 18080
rect 5582 17926 5634 17978
rect 5646 17926 5698 17978
rect 5710 17926 5762 17978
rect 5774 17926 5826 17978
rect 5838 17926 5890 17978
rect 14846 17926 14898 17978
rect 14910 17926 14962 17978
rect 14974 17926 15026 17978
rect 15038 17926 15090 17978
rect 15102 17926 15154 17978
rect 24110 17926 24162 17978
rect 24174 17926 24226 17978
rect 24238 17926 24290 17978
rect 24302 17926 24354 17978
rect 24366 17926 24418 17978
rect 8116 17867 8168 17876
rect 8116 17833 8125 17867
rect 8125 17833 8159 17867
rect 8159 17833 8168 17867
rect 8116 17824 8168 17833
rect 10600 17867 10652 17876
rect 10600 17833 10609 17867
rect 10609 17833 10643 17867
rect 10643 17833 10652 17867
rect 10600 17824 10652 17833
rect 11152 17867 11204 17876
rect 11152 17833 11161 17867
rect 11161 17833 11195 17867
rect 11195 17833 11204 17867
rect 11152 17824 11204 17833
rect 12716 17824 12768 17876
rect 13360 17824 13412 17876
rect 17592 17824 17644 17876
rect 10324 17799 10376 17808
rect 10324 17765 10333 17799
rect 10333 17765 10367 17799
rect 10367 17765 10376 17799
rect 10324 17756 10376 17765
rect 12992 17799 13044 17808
rect 12992 17765 13001 17799
rect 13001 17765 13035 17799
rect 13035 17765 13044 17799
rect 12992 17756 13044 17765
rect 18144 17824 18196 17876
rect 18604 17824 18656 17876
rect 21640 17824 21692 17876
rect 23020 17824 23072 17876
rect 15476 17731 15528 17740
rect 6000 17663 6052 17672
rect 6000 17629 6009 17663
rect 6009 17629 6043 17663
rect 6043 17629 6052 17663
rect 6000 17620 6052 17629
rect 9036 17620 9088 17672
rect 10968 17663 11020 17672
rect 10968 17629 10977 17663
rect 10977 17629 11011 17663
rect 11011 17629 11020 17663
rect 10968 17620 11020 17629
rect 11980 17620 12032 17672
rect 12808 17620 12860 17672
rect 6092 17552 6144 17604
rect 8024 17595 8076 17604
rect 8024 17561 8033 17595
rect 8033 17561 8067 17595
rect 8067 17561 8076 17595
rect 8024 17552 8076 17561
rect 8668 17552 8720 17604
rect 12624 17595 12676 17604
rect 12624 17561 12633 17595
rect 12633 17561 12667 17595
rect 12667 17561 12676 17595
rect 12624 17552 12676 17561
rect 14188 17620 14240 17672
rect 14461 17657 14513 17666
rect 14461 17623 14470 17657
rect 14470 17623 14504 17657
rect 14504 17623 14513 17657
rect 14461 17614 14513 17623
rect 14648 17620 14700 17672
rect 7380 17527 7432 17536
rect 7380 17493 7389 17527
rect 7389 17493 7423 17527
rect 7423 17493 7432 17527
rect 7380 17484 7432 17493
rect 12440 17484 12492 17536
rect 13544 17552 13596 17604
rect 15476 17697 15485 17731
rect 15485 17697 15519 17731
rect 15519 17697 15528 17731
rect 15476 17688 15528 17697
rect 15200 17620 15252 17672
rect 15660 17663 15712 17672
rect 15660 17629 15668 17663
rect 15668 17629 15702 17663
rect 15702 17629 15712 17663
rect 15660 17620 15712 17629
rect 19340 17688 19392 17740
rect 19984 17688 20036 17740
rect 20352 17688 20404 17740
rect 16488 17552 16540 17604
rect 18512 17552 18564 17604
rect 18604 17595 18656 17604
rect 18604 17561 18613 17595
rect 18613 17561 18647 17595
rect 18647 17561 18656 17595
rect 18604 17552 18656 17561
rect 19892 17620 19944 17672
rect 20628 17756 20680 17808
rect 20720 17756 20772 17808
rect 22284 17799 22336 17808
rect 22284 17765 22293 17799
rect 22293 17765 22327 17799
rect 22327 17765 22336 17799
rect 22284 17756 22336 17765
rect 22744 17688 22796 17740
rect 20904 17663 20956 17672
rect 20904 17629 20913 17663
rect 20913 17629 20947 17663
rect 20947 17629 20956 17663
rect 20904 17620 20956 17629
rect 21272 17620 21324 17672
rect 23112 17663 23164 17672
rect 23112 17629 23121 17663
rect 23121 17629 23155 17663
rect 23155 17629 23164 17663
rect 23112 17620 23164 17629
rect 14096 17527 14148 17536
rect 14096 17493 14105 17527
rect 14105 17493 14139 17527
rect 14139 17493 14148 17527
rect 14096 17484 14148 17493
rect 14648 17484 14700 17536
rect 16120 17484 16172 17536
rect 16304 17484 16356 17536
rect 18236 17484 18288 17536
rect 20260 17527 20312 17536
rect 20260 17493 20269 17527
rect 20269 17493 20303 17527
rect 20303 17493 20312 17527
rect 20260 17484 20312 17493
rect 21732 17552 21784 17604
rect 22468 17595 22520 17604
rect 22468 17561 22477 17595
rect 22477 17561 22511 17595
rect 22511 17561 22520 17595
rect 22468 17552 22520 17561
rect 21916 17484 21968 17536
rect 23020 17552 23072 17604
rect 23848 17552 23900 17604
rect 23204 17484 23256 17536
rect 23388 17484 23440 17536
rect 25412 17484 25464 17536
rect 10214 17382 10266 17434
rect 10278 17382 10330 17434
rect 10342 17382 10394 17434
rect 10406 17382 10458 17434
rect 10470 17382 10522 17434
rect 19478 17382 19530 17434
rect 19542 17382 19594 17434
rect 19606 17382 19658 17434
rect 19670 17382 19722 17434
rect 19734 17382 19786 17434
rect 6092 17280 6144 17332
rect 8668 17323 8720 17332
rect 8668 17289 8677 17323
rect 8677 17289 8711 17323
rect 8711 17289 8720 17323
rect 8668 17280 8720 17289
rect 9864 17323 9916 17332
rect 9864 17289 9873 17323
rect 9873 17289 9907 17323
rect 9907 17289 9916 17323
rect 9864 17280 9916 17289
rect 7380 17255 7432 17264
rect 7380 17221 7389 17255
rect 7389 17221 7423 17255
rect 7423 17221 7432 17255
rect 7380 17212 7432 17221
rect 9128 17187 9180 17196
rect 9128 17153 9137 17187
rect 9137 17153 9171 17187
rect 9171 17153 9180 17187
rect 9128 17144 9180 17153
rect 6644 17076 6696 17128
rect 7472 17119 7524 17128
rect 7472 17085 7481 17119
rect 7481 17085 7515 17119
rect 7515 17085 7524 17119
rect 7472 17076 7524 17085
rect 7840 17076 7892 17128
rect 8024 17076 8076 17128
rect 9312 17119 9364 17128
rect 9312 17085 9321 17119
rect 9321 17085 9355 17119
rect 9355 17085 9364 17119
rect 9312 17076 9364 17085
rect 10600 17212 10652 17264
rect 10968 17212 11020 17264
rect 13268 17280 13320 17332
rect 15568 17280 15620 17332
rect 18236 17280 18288 17332
rect 18512 17280 18564 17332
rect 21088 17280 21140 17332
rect 23020 17280 23072 17332
rect 25412 17280 25464 17332
rect 11612 17212 11664 17264
rect 12348 17212 12400 17264
rect 12256 17144 12308 17196
rect 14004 17144 14056 17196
rect 14464 17187 14516 17196
rect 11060 17076 11112 17128
rect 11520 17119 11572 17128
rect 11520 17085 11529 17119
rect 11529 17085 11563 17119
rect 11563 17085 11572 17119
rect 11520 17076 11572 17085
rect 13636 17076 13688 17128
rect 1400 17051 1452 17060
rect 1400 17017 1409 17051
rect 1409 17017 1443 17051
rect 1443 17017 1452 17051
rect 1400 17008 1452 17017
rect 10324 16983 10376 16992
rect 10324 16949 10333 16983
rect 10333 16949 10367 16983
rect 10367 16949 10376 16983
rect 10324 16940 10376 16949
rect 12992 17008 13044 17060
rect 14464 17153 14473 17187
rect 14473 17153 14507 17187
rect 14507 17153 14516 17187
rect 14464 17144 14516 17153
rect 15752 17144 15804 17196
rect 14556 17076 14608 17128
rect 15476 17076 15528 17128
rect 16120 17144 16172 17196
rect 17592 17187 17644 17196
rect 17224 17076 17276 17128
rect 17592 17153 17601 17187
rect 17601 17153 17635 17187
rect 17635 17153 17644 17187
rect 17592 17144 17644 17153
rect 17960 17144 18012 17196
rect 20260 17212 20312 17264
rect 18696 17144 18748 17196
rect 19340 17144 19392 17196
rect 21180 17144 21232 17196
rect 21364 17144 21416 17196
rect 22192 17187 22244 17196
rect 22192 17153 22201 17187
rect 22201 17153 22235 17187
rect 22235 17153 22244 17187
rect 22192 17144 22244 17153
rect 23204 17187 23256 17196
rect 23204 17153 23213 17187
rect 23213 17153 23247 17187
rect 23247 17153 23256 17187
rect 23204 17144 23256 17153
rect 23848 17144 23900 17196
rect 28356 17187 28408 17196
rect 28356 17153 28365 17187
rect 28365 17153 28399 17187
rect 28399 17153 28408 17187
rect 28356 17144 28408 17153
rect 23020 17076 23072 17128
rect 23756 17076 23808 17128
rect 23940 17119 23992 17128
rect 23940 17085 23949 17119
rect 23949 17085 23983 17119
rect 23983 17085 23992 17119
rect 23940 17076 23992 17085
rect 11888 16940 11940 16992
rect 13268 16940 13320 16992
rect 13820 16983 13872 16992
rect 13820 16949 13829 16983
rect 13829 16949 13863 16983
rect 13863 16949 13872 16983
rect 13820 16940 13872 16949
rect 19616 17008 19668 17060
rect 14464 16940 14516 16992
rect 15200 16940 15252 16992
rect 17500 16940 17552 16992
rect 19064 16983 19116 16992
rect 19064 16949 19073 16983
rect 19073 16949 19107 16983
rect 19107 16949 19116 16983
rect 19064 16940 19116 16949
rect 19524 16940 19576 16992
rect 20352 16940 20404 16992
rect 20720 16940 20772 16992
rect 21732 16940 21784 16992
rect 21916 16940 21968 16992
rect 5582 16838 5634 16890
rect 5646 16838 5698 16890
rect 5710 16838 5762 16890
rect 5774 16838 5826 16890
rect 5838 16838 5890 16890
rect 14846 16838 14898 16890
rect 14910 16838 14962 16890
rect 14974 16838 15026 16890
rect 15038 16838 15090 16890
rect 15102 16838 15154 16890
rect 24110 16838 24162 16890
rect 24174 16838 24226 16890
rect 24238 16838 24290 16890
rect 24302 16838 24354 16890
rect 24366 16838 24418 16890
rect 7472 16736 7524 16788
rect 7656 16736 7708 16788
rect 9036 16600 9088 16652
rect 9864 16736 9916 16788
rect 10692 16736 10744 16788
rect 10876 16736 10928 16788
rect 11060 16736 11112 16788
rect 12164 16779 12216 16788
rect 12164 16745 12173 16779
rect 12173 16745 12207 16779
rect 12207 16745 12216 16779
rect 12164 16736 12216 16745
rect 15844 16736 15896 16788
rect 16856 16779 16908 16788
rect 16856 16745 16865 16779
rect 16865 16745 16899 16779
rect 16899 16745 16908 16779
rect 16856 16736 16908 16745
rect 17224 16779 17276 16788
rect 17224 16745 17233 16779
rect 17233 16745 17267 16779
rect 17267 16745 17276 16779
rect 17224 16736 17276 16745
rect 18328 16736 18380 16788
rect 19248 16736 19300 16788
rect 19524 16779 19576 16788
rect 19524 16745 19533 16779
rect 19533 16745 19567 16779
rect 19567 16745 19576 16779
rect 19524 16736 19576 16745
rect 19616 16736 19668 16788
rect 23848 16779 23900 16788
rect 23848 16745 23857 16779
rect 23857 16745 23891 16779
rect 23891 16745 23900 16779
rect 23848 16736 23900 16745
rect 25044 16779 25096 16788
rect 25044 16745 25053 16779
rect 25053 16745 25087 16779
rect 25087 16745 25096 16779
rect 25044 16736 25096 16745
rect 13636 16668 13688 16720
rect 10324 16600 10376 16652
rect 4620 16532 4672 16584
rect 9312 16532 9364 16584
rect 9772 16532 9824 16584
rect 13912 16600 13964 16652
rect 8300 16507 8352 16516
rect 8300 16473 8318 16507
rect 8318 16473 8352 16507
rect 8300 16464 8352 16473
rect 10784 16532 10836 16584
rect 10876 16464 10928 16516
rect 11152 16464 11204 16516
rect 11888 16507 11940 16516
rect 11888 16473 11897 16507
rect 11897 16473 11931 16507
rect 11931 16473 11940 16507
rect 11888 16464 11940 16473
rect 13360 16575 13412 16584
rect 13360 16541 13369 16575
rect 13369 16541 13403 16575
rect 13403 16541 13412 16575
rect 13360 16532 13412 16541
rect 13544 16575 13596 16584
rect 13544 16541 13553 16575
rect 13553 16541 13587 16575
rect 13587 16541 13596 16575
rect 13544 16532 13596 16541
rect 14096 16532 14148 16584
rect 15016 16668 15068 16720
rect 14556 16643 14608 16652
rect 14556 16609 14565 16643
rect 14565 16609 14599 16643
rect 14599 16609 14608 16643
rect 14556 16600 14608 16609
rect 15752 16643 15804 16652
rect 15752 16609 15761 16643
rect 15761 16609 15795 16643
rect 15795 16609 15804 16643
rect 15752 16600 15804 16609
rect 14372 16575 14424 16584
rect 14372 16541 14381 16575
rect 14381 16541 14415 16575
rect 14415 16541 14424 16575
rect 14648 16575 14700 16584
rect 14372 16532 14424 16541
rect 14648 16541 14657 16575
rect 14657 16541 14691 16575
rect 14691 16541 14700 16575
rect 14648 16532 14700 16541
rect 15108 16575 15160 16584
rect 15108 16541 15117 16575
rect 15117 16541 15151 16575
rect 15151 16541 15160 16575
rect 15108 16532 15160 16541
rect 15476 16532 15528 16584
rect 15660 16575 15712 16584
rect 15660 16541 15669 16575
rect 15669 16541 15703 16575
rect 15703 16541 15712 16575
rect 15660 16532 15712 16541
rect 15936 16575 15988 16584
rect 15936 16541 15945 16575
rect 15945 16541 15979 16575
rect 15979 16541 15988 16575
rect 15936 16532 15988 16541
rect 22652 16711 22704 16720
rect 17316 16600 17368 16652
rect 1492 16439 1544 16448
rect 1492 16405 1501 16439
rect 1501 16405 1535 16439
rect 1535 16405 1544 16439
rect 1492 16396 1544 16405
rect 9220 16439 9272 16448
rect 9220 16405 9229 16439
rect 9229 16405 9263 16439
rect 9263 16405 9272 16439
rect 9220 16396 9272 16405
rect 10692 16396 10744 16448
rect 12900 16439 12952 16448
rect 12900 16405 12909 16439
rect 12909 16405 12943 16439
rect 12943 16405 12952 16439
rect 12900 16396 12952 16405
rect 16304 16464 16356 16516
rect 16764 16507 16816 16516
rect 16764 16473 16773 16507
rect 16773 16473 16807 16507
rect 16807 16473 16816 16507
rect 16764 16464 16816 16473
rect 17224 16532 17276 16584
rect 20260 16600 20312 16652
rect 22652 16677 22661 16711
rect 22661 16677 22695 16711
rect 22695 16677 22704 16711
rect 22652 16668 22704 16677
rect 19248 16575 19300 16584
rect 18420 16464 18472 16516
rect 13544 16396 13596 16448
rect 15108 16396 15160 16448
rect 15200 16396 15252 16448
rect 16396 16396 16448 16448
rect 17776 16396 17828 16448
rect 18052 16396 18104 16448
rect 18236 16396 18288 16448
rect 18696 16396 18748 16448
rect 19248 16541 19257 16575
rect 19257 16541 19291 16575
rect 19291 16541 19300 16575
rect 19248 16532 19300 16541
rect 19064 16464 19116 16516
rect 20168 16532 20220 16584
rect 21088 16532 21140 16584
rect 21732 16575 21784 16584
rect 21732 16541 21741 16575
rect 21741 16541 21775 16575
rect 21775 16541 21784 16575
rect 21732 16532 21784 16541
rect 21916 16575 21968 16584
rect 21916 16541 21925 16575
rect 21925 16541 21959 16575
rect 21959 16541 21968 16575
rect 21916 16532 21968 16541
rect 23296 16600 23348 16652
rect 28356 16643 28408 16652
rect 28356 16609 28365 16643
rect 28365 16609 28399 16643
rect 28399 16609 28408 16643
rect 28356 16600 28408 16609
rect 22468 16532 22520 16584
rect 23020 16532 23072 16584
rect 23388 16575 23440 16584
rect 23388 16541 23397 16575
rect 23397 16541 23431 16575
rect 23431 16541 23440 16575
rect 23388 16532 23440 16541
rect 20720 16507 20772 16516
rect 20720 16473 20729 16507
rect 20729 16473 20763 16507
rect 20763 16473 20772 16507
rect 20720 16464 20772 16473
rect 21180 16507 21232 16516
rect 21180 16473 21189 16507
rect 21189 16473 21223 16507
rect 21223 16473 21232 16507
rect 21180 16464 21232 16473
rect 22192 16464 22244 16516
rect 22560 16464 22612 16516
rect 23112 16464 23164 16516
rect 23572 16575 23624 16584
rect 23572 16541 23581 16575
rect 23581 16541 23615 16575
rect 23615 16541 23624 16575
rect 23572 16532 23624 16541
rect 25044 16532 25096 16584
rect 23756 16464 23808 16516
rect 24584 16507 24636 16516
rect 24584 16473 24593 16507
rect 24593 16473 24627 16507
rect 24627 16473 24636 16507
rect 24584 16464 24636 16473
rect 19892 16396 19944 16448
rect 21088 16396 21140 16448
rect 23664 16396 23716 16448
rect 10214 16294 10266 16346
rect 10278 16294 10330 16346
rect 10342 16294 10394 16346
rect 10406 16294 10458 16346
rect 10470 16294 10522 16346
rect 19478 16294 19530 16346
rect 19542 16294 19594 16346
rect 19606 16294 19658 16346
rect 19670 16294 19722 16346
rect 19734 16294 19786 16346
rect 7656 16235 7708 16244
rect 7656 16201 7665 16235
rect 7665 16201 7699 16235
rect 7699 16201 7708 16235
rect 7656 16192 7708 16201
rect 9312 16192 9364 16244
rect 11888 16192 11940 16244
rect 11980 16192 12032 16244
rect 5908 16056 5960 16108
rect 6644 16099 6696 16108
rect 6644 16065 6653 16099
rect 6653 16065 6687 16099
rect 6687 16065 6696 16099
rect 6644 16056 6696 16065
rect 9772 16124 9824 16176
rect 9220 16056 9272 16108
rect 9588 16099 9640 16108
rect 9588 16065 9622 16099
rect 9622 16065 9640 16099
rect 9588 16056 9640 16065
rect 11244 16056 11296 16108
rect 11428 16056 11480 16108
rect 11704 16056 11756 16108
rect 13268 16167 13320 16176
rect 13268 16133 13277 16167
rect 13277 16133 13311 16167
rect 13311 16133 13320 16167
rect 13268 16124 13320 16133
rect 13544 16124 13596 16176
rect 7656 15920 7708 15972
rect 7840 16031 7892 16040
rect 7840 15997 7849 16031
rect 7849 15997 7883 16031
rect 7883 15997 7892 16031
rect 9312 16031 9364 16040
rect 7840 15988 7892 15997
rect 9312 15997 9321 16031
rect 9321 15997 9355 16031
rect 9355 15997 9364 16031
rect 9312 15988 9364 15997
rect 5172 15852 5224 15904
rect 8484 15852 8536 15904
rect 9036 15895 9088 15904
rect 9036 15861 9045 15895
rect 9045 15861 9079 15895
rect 9079 15861 9088 15895
rect 9036 15852 9088 15861
rect 11152 15920 11204 15972
rect 12256 15988 12308 16040
rect 13912 16124 13964 16176
rect 14004 16099 14056 16108
rect 14004 16065 14013 16099
rect 14013 16065 14047 16099
rect 14047 16065 14056 16099
rect 14004 16056 14056 16065
rect 15476 16192 15528 16244
rect 14464 16124 14516 16176
rect 16948 16192 17000 16244
rect 14556 16099 14608 16108
rect 14556 16065 14565 16099
rect 14565 16065 14599 16099
rect 14599 16065 14608 16099
rect 14556 16056 14608 16065
rect 16672 16124 16724 16176
rect 15108 16099 15160 16108
rect 15108 16065 15117 16099
rect 15117 16065 15151 16099
rect 15151 16065 15160 16099
rect 15108 16056 15160 16065
rect 15200 16099 15252 16108
rect 15200 16065 15209 16099
rect 15209 16065 15243 16099
rect 15243 16065 15252 16099
rect 16028 16099 16080 16108
rect 15200 16056 15252 16065
rect 16028 16065 16037 16099
rect 16037 16065 16071 16099
rect 16071 16065 16080 16099
rect 16028 16056 16080 16065
rect 16488 16056 16540 16108
rect 17776 16192 17828 16244
rect 19156 16192 19208 16244
rect 19340 16192 19392 16244
rect 21180 16192 21232 16244
rect 24584 16192 24636 16244
rect 17316 16124 17368 16176
rect 17868 16099 17920 16108
rect 15752 15988 15804 16040
rect 16120 16031 16172 16040
rect 15016 15920 15068 15972
rect 15384 15963 15436 15972
rect 15384 15929 15393 15963
rect 15393 15929 15427 15963
rect 15427 15929 15436 15963
rect 15384 15920 15436 15929
rect 16120 15997 16129 16031
rect 16129 15997 16163 16031
rect 16163 15997 16172 16031
rect 16120 15988 16172 15997
rect 16856 15988 16908 16040
rect 17868 16065 17877 16099
rect 17877 16065 17911 16099
rect 17911 16065 17920 16099
rect 17868 16056 17920 16065
rect 18328 16099 18380 16108
rect 18328 16065 18337 16099
rect 18337 16065 18371 16099
rect 18371 16065 18380 16099
rect 18328 16056 18380 16065
rect 18788 16056 18840 16108
rect 19156 16056 19208 16108
rect 19892 16056 19944 16108
rect 20076 16099 20128 16108
rect 20076 16065 20085 16099
rect 20085 16065 20119 16099
rect 20119 16065 20128 16099
rect 20076 16056 20128 16065
rect 10692 15895 10744 15904
rect 10692 15861 10701 15895
rect 10701 15861 10735 15895
rect 10735 15861 10744 15895
rect 10692 15852 10744 15861
rect 10876 15852 10928 15904
rect 11244 15852 11296 15904
rect 12808 15895 12860 15904
rect 12808 15861 12817 15895
rect 12817 15861 12851 15895
rect 12851 15861 12860 15895
rect 12808 15852 12860 15861
rect 13544 15852 13596 15904
rect 17776 15852 17828 15904
rect 20352 15988 20404 16040
rect 21088 16099 21140 16108
rect 21088 16065 21097 16099
rect 21097 16065 21131 16099
rect 21131 16065 21140 16099
rect 21088 16056 21140 16065
rect 21732 16056 21784 16108
rect 22008 16099 22060 16108
rect 22008 16065 22017 16099
rect 22017 16065 22051 16099
rect 22051 16065 22060 16099
rect 22008 16056 22060 16065
rect 22468 16124 22520 16176
rect 23020 16099 23072 16108
rect 23020 16065 23029 16099
rect 23029 16065 23063 16099
rect 23063 16065 23072 16099
rect 23020 16056 23072 16065
rect 23204 16099 23256 16108
rect 23204 16065 23208 16099
rect 23208 16065 23242 16099
rect 23242 16065 23256 16099
rect 23204 16056 23256 16065
rect 19432 15963 19484 15972
rect 19432 15929 19441 15963
rect 19441 15929 19475 15963
rect 19475 15929 19484 15963
rect 19432 15920 19484 15929
rect 20996 15920 21048 15972
rect 21088 15920 21140 15972
rect 22100 15920 22152 15972
rect 23112 15920 23164 15972
rect 23388 16099 23440 16108
rect 23388 16065 23397 16099
rect 23397 16065 23431 16099
rect 23431 16065 23440 16099
rect 23388 16056 23440 16065
rect 26424 16056 26476 16108
rect 23940 16031 23992 16040
rect 23940 15997 23949 16031
rect 23949 15997 23983 16031
rect 23983 15997 23992 16031
rect 23940 15988 23992 15997
rect 19892 15852 19944 15904
rect 21548 15852 21600 15904
rect 22836 15852 22888 15904
rect 5582 15750 5634 15802
rect 5646 15750 5698 15802
rect 5710 15750 5762 15802
rect 5774 15750 5826 15802
rect 5838 15750 5890 15802
rect 14846 15750 14898 15802
rect 14910 15750 14962 15802
rect 14974 15750 15026 15802
rect 15038 15750 15090 15802
rect 15102 15750 15154 15802
rect 24110 15750 24162 15802
rect 24174 15750 24226 15802
rect 24238 15750 24290 15802
rect 24302 15750 24354 15802
rect 24366 15750 24418 15802
rect 5908 15648 5960 15700
rect 8300 15691 8352 15700
rect 8300 15657 8309 15691
rect 8309 15657 8343 15691
rect 8343 15657 8352 15691
rect 8300 15648 8352 15657
rect 9588 15648 9640 15700
rect 11704 15691 11756 15700
rect 11704 15657 11713 15691
rect 11713 15657 11747 15691
rect 11747 15657 11756 15691
rect 11704 15648 11756 15657
rect 11888 15648 11940 15700
rect 13544 15691 13596 15700
rect 7656 15580 7708 15632
rect 7288 15512 7340 15564
rect 7840 15555 7892 15564
rect 7840 15521 7849 15555
rect 7849 15521 7883 15555
rect 7883 15521 7892 15555
rect 7840 15512 7892 15521
rect 10876 15512 10928 15564
rect 13544 15657 13553 15691
rect 13553 15657 13587 15691
rect 13587 15657 13596 15691
rect 13544 15648 13596 15657
rect 15200 15648 15252 15700
rect 22008 15648 22060 15700
rect 22192 15648 22244 15700
rect 22928 15648 22980 15700
rect 20536 15623 20588 15632
rect 20536 15589 20545 15623
rect 20545 15589 20579 15623
rect 20579 15589 20588 15623
rect 20536 15580 20588 15589
rect 22468 15580 22520 15632
rect 23020 15580 23072 15632
rect 23204 15580 23256 15632
rect 17868 15555 17920 15564
rect 17868 15521 17877 15555
rect 17877 15521 17911 15555
rect 17911 15521 17920 15555
rect 17868 15512 17920 15521
rect 19432 15512 19484 15564
rect 20352 15555 20404 15564
rect 20352 15521 20361 15555
rect 20361 15521 20395 15555
rect 20395 15521 20404 15555
rect 21456 15555 21508 15564
rect 20352 15512 20404 15521
rect 21456 15521 21465 15555
rect 21465 15521 21499 15555
rect 21499 15521 21508 15555
rect 21456 15512 21508 15521
rect 5172 15487 5224 15496
rect 5172 15453 5181 15487
rect 5181 15453 5215 15487
rect 5215 15453 5224 15487
rect 5172 15444 5224 15453
rect 5632 15487 5684 15496
rect 5632 15453 5641 15487
rect 5641 15453 5675 15487
rect 5675 15453 5684 15487
rect 5632 15444 5684 15453
rect 7656 15487 7708 15496
rect 7656 15453 7665 15487
rect 7665 15453 7699 15487
rect 7699 15453 7708 15487
rect 7656 15444 7708 15453
rect 7748 15487 7800 15496
rect 7748 15453 7757 15487
rect 7757 15453 7791 15487
rect 7791 15453 7800 15487
rect 8484 15487 8536 15496
rect 7748 15444 7800 15453
rect 8484 15453 8493 15487
rect 8493 15453 8527 15487
rect 8527 15453 8536 15487
rect 8484 15444 8536 15453
rect 9036 15444 9088 15496
rect 11244 15487 11296 15496
rect 11244 15453 11253 15487
rect 11253 15453 11287 15487
rect 11287 15453 11296 15487
rect 11244 15444 11296 15453
rect 15844 15487 15896 15496
rect 7196 15376 7248 15428
rect 12348 15376 12400 15428
rect 12532 15376 12584 15428
rect 15844 15453 15853 15487
rect 15853 15453 15887 15487
rect 15887 15453 15896 15487
rect 15844 15444 15896 15453
rect 16028 15444 16080 15496
rect 18420 15444 18472 15496
rect 20076 15444 20128 15496
rect 21088 15444 21140 15496
rect 22376 15487 22428 15496
rect 22376 15453 22385 15487
rect 22385 15453 22419 15487
rect 22419 15453 22428 15487
rect 22376 15444 22428 15453
rect 22652 15444 22704 15496
rect 23848 15648 23900 15700
rect 28172 15648 28224 15700
rect 23940 15512 23992 15564
rect 25136 15444 25188 15496
rect 28356 15487 28408 15496
rect 28356 15453 28365 15487
rect 28365 15453 28399 15487
rect 28399 15453 28408 15487
rect 28356 15444 28408 15453
rect 10692 15308 10744 15360
rect 13636 15376 13688 15428
rect 15016 15376 15068 15428
rect 20720 15376 20772 15428
rect 21916 15419 21968 15428
rect 14096 15308 14148 15360
rect 14648 15308 14700 15360
rect 15384 15308 15436 15360
rect 17132 15351 17184 15360
rect 17132 15317 17141 15351
rect 17141 15317 17175 15351
rect 17175 15317 17184 15351
rect 17132 15308 17184 15317
rect 21916 15385 21925 15419
rect 21925 15385 21959 15419
rect 21959 15385 21968 15419
rect 21916 15376 21968 15385
rect 22560 15308 22612 15360
rect 22928 15308 22980 15360
rect 23572 15376 23624 15428
rect 23940 15308 23992 15360
rect 10214 15206 10266 15258
rect 10278 15206 10330 15258
rect 10342 15206 10394 15258
rect 10406 15206 10458 15258
rect 10470 15206 10522 15258
rect 19478 15206 19530 15258
rect 19542 15206 19594 15258
rect 19606 15206 19658 15258
rect 19670 15206 19722 15258
rect 19734 15206 19786 15258
rect 11152 15104 11204 15156
rect 12532 15147 12584 15156
rect 12532 15113 12541 15147
rect 12541 15113 12575 15147
rect 12575 15113 12584 15147
rect 12532 15104 12584 15113
rect 15016 15147 15068 15156
rect 15016 15113 15025 15147
rect 15025 15113 15059 15147
rect 15059 15113 15068 15147
rect 15016 15104 15068 15113
rect 8208 15036 8260 15088
rect 10600 15036 10652 15088
rect 15568 15036 15620 15088
rect 5632 14968 5684 15020
rect 6000 14968 6052 15020
rect 8116 15011 8168 15020
rect 8116 14977 8150 15011
rect 8150 14977 8168 15011
rect 8116 14968 8168 14977
rect 9312 14968 9364 15020
rect 11428 14968 11480 15020
rect 11980 14968 12032 15020
rect 12348 15011 12400 15020
rect 12348 14977 12357 15011
rect 12357 14977 12391 15011
rect 12391 14977 12400 15011
rect 12348 14968 12400 14977
rect 13544 15011 13596 15020
rect 13544 14977 13553 15011
rect 13553 14977 13587 15011
rect 13587 14977 13596 15011
rect 13544 14968 13596 14977
rect 13636 14900 13688 14952
rect 13912 14968 13964 15020
rect 14280 14968 14332 15020
rect 15200 14968 15252 15020
rect 15476 15011 15528 15020
rect 15476 14977 15485 15011
rect 15485 14977 15519 15011
rect 15519 14977 15528 15011
rect 16212 15104 16264 15156
rect 16764 15104 16816 15156
rect 17776 15147 17828 15156
rect 17776 15113 17785 15147
rect 17785 15113 17819 15147
rect 17819 15113 17828 15147
rect 17776 15104 17828 15113
rect 16028 15036 16080 15088
rect 15476 14968 15528 14977
rect 15752 14900 15804 14952
rect 12900 14832 12952 14884
rect 9404 14764 9456 14816
rect 11336 14764 11388 14816
rect 13268 14807 13320 14816
rect 13268 14773 13277 14807
rect 13277 14773 13311 14807
rect 13311 14773 13320 14807
rect 13268 14764 13320 14773
rect 14188 14764 14240 14816
rect 14464 14832 14516 14884
rect 15844 14832 15896 14884
rect 16212 14968 16264 15020
rect 16488 14968 16540 15020
rect 16856 14968 16908 15020
rect 16396 14900 16448 14952
rect 19800 15036 19852 15088
rect 20444 15104 20496 15156
rect 21272 15147 21324 15156
rect 21272 15113 21281 15147
rect 21281 15113 21315 15147
rect 21315 15113 21324 15147
rect 21272 15104 21324 15113
rect 22008 15147 22060 15156
rect 22008 15113 22017 15147
rect 22017 15113 22051 15147
rect 22051 15113 22060 15147
rect 22008 15104 22060 15113
rect 25136 15147 25188 15156
rect 25136 15113 25145 15147
rect 25145 15113 25179 15147
rect 25179 15113 25188 15147
rect 25136 15104 25188 15113
rect 19340 14968 19392 15020
rect 18328 14900 18380 14952
rect 20628 15036 20680 15088
rect 21916 15036 21968 15088
rect 23940 15036 23992 15088
rect 24860 15079 24912 15088
rect 24860 15045 24869 15079
rect 24869 15045 24903 15079
rect 24903 15045 24912 15079
rect 24860 15036 24912 15045
rect 20720 15011 20772 15020
rect 20720 14977 20729 15011
rect 20729 14977 20763 15011
rect 20763 14977 20772 15011
rect 20720 14968 20772 14977
rect 20996 14968 21048 15020
rect 21180 14968 21232 15020
rect 21732 14968 21784 15020
rect 23020 14968 23072 15020
rect 23756 15011 23808 15020
rect 20536 14943 20588 14952
rect 20536 14909 20545 14943
rect 20545 14909 20579 14943
rect 20579 14909 20588 14943
rect 20536 14900 20588 14909
rect 22008 14900 22060 14952
rect 22928 14900 22980 14952
rect 23756 14977 23765 15011
rect 23765 14977 23799 15011
rect 23799 14977 23808 15011
rect 23756 14968 23808 14977
rect 23572 14900 23624 14952
rect 18788 14832 18840 14884
rect 19064 14832 19116 14884
rect 17684 14764 17736 14816
rect 18052 14764 18104 14816
rect 18512 14807 18564 14816
rect 18512 14773 18521 14807
rect 18521 14773 18555 14807
rect 18555 14773 18564 14807
rect 18512 14764 18564 14773
rect 18972 14764 19024 14816
rect 21088 14832 21140 14884
rect 21180 14832 21232 14884
rect 24032 14807 24084 14816
rect 24032 14773 24041 14807
rect 24041 14773 24075 14807
rect 24075 14773 24084 14807
rect 24032 14764 24084 14773
rect 5582 14662 5634 14714
rect 5646 14662 5698 14714
rect 5710 14662 5762 14714
rect 5774 14662 5826 14714
rect 5838 14662 5890 14714
rect 14846 14662 14898 14714
rect 14910 14662 14962 14714
rect 14974 14662 15026 14714
rect 15038 14662 15090 14714
rect 15102 14662 15154 14714
rect 24110 14662 24162 14714
rect 24174 14662 24226 14714
rect 24238 14662 24290 14714
rect 24302 14662 24354 14714
rect 24366 14662 24418 14714
rect 11980 14560 12032 14612
rect 12900 14560 12952 14612
rect 13084 14603 13136 14612
rect 13084 14569 13093 14603
rect 13093 14569 13127 14603
rect 13127 14569 13136 14603
rect 13084 14560 13136 14569
rect 8668 14492 8720 14544
rect 12624 14492 12676 14544
rect 13544 14492 13596 14544
rect 15476 14560 15528 14612
rect 15568 14560 15620 14612
rect 15660 14492 15712 14544
rect 16764 14560 16816 14612
rect 18052 14560 18104 14612
rect 18880 14560 18932 14612
rect 19524 14560 19576 14612
rect 19984 14560 20036 14612
rect 21364 14603 21416 14612
rect 21364 14569 21373 14603
rect 21373 14569 21407 14603
rect 21407 14569 21416 14603
rect 21364 14560 21416 14569
rect 22560 14603 22612 14612
rect 22560 14569 22569 14603
rect 22569 14569 22603 14603
rect 22603 14569 22612 14603
rect 22560 14560 22612 14569
rect 23112 14560 23164 14612
rect 23480 14560 23532 14612
rect 26056 14560 26108 14612
rect 16396 14492 16448 14544
rect 16488 14492 16540 14544
rect 17776 14492 17828 14544
rect 18604 14492 18656 14544
rect 18788 14535 18840 14544
rect 18788 14501 18797 14535
rect 18797 14501 18831 14535
rect 18831 14501 18840 14535
rect 18788 14492 18840 14501
rect 4436 14356 4488 14408
rect 8300 14356 8352 14408
rect 9404 14356 9456 14408
rect 11980 14356 12032 14408
rect 6920 14288 6972 14340
rect 14188 14424 14240 14476
rect 8484 14220 8536 14272
rect 9496 14263 9548 14272
rect 9496 14229 9505 14263
rect 9505 14229 9539 14263
rect 9539 14229 9548 14263
rect 9496 14220 9548 14229
rect 14280 14356 14332 14408
rect 15476 14424 15528 14476
rect 16028 14424 16080 14476
rect 16120 14467 16172 14476
rect 16120 14433 16129 14467
rect 16129 14433 16163 14467
rect 16163 14433 16172 14467
rect 16120 14424 16172 14433
rect 14648 14356 14700 14408
rect 15384 14356 15436 14408
rect 18328 14424 18380 14476
rect 19340 14467 19392 14476
rect 19340 14433 19349 14467
rect 19349 14433 19383 14467
rect 19383 14433 19392 14467
rect 19340 14424 19392 14433
rect 20536 14492 20588 14544
rect 20628 14492 20680 14544
rect 24032 14492 24084 14544
rect 21456 14424 21508 14476
rect 16948 14399 17000 14408
rect 15200 14288 15252 14340
rect 13912 14220 13964 14272
rect 14280 14220 14332 14272
rect 14464 14220 14516 14272
rect 14648 14220 14700 14272
rect 15936 14288 15988 14340
rect 16396 14288 16448 14340
rect 16948 14365 16957 14399
rect 16957 14365 16991 14399
rect 16991 14365 17000 14399
rect 16948 14356 17000 14365
rect 17040 14399 17092 14408
rect 17040 14365 17049 14399
rect 17049 14365 17083 14399
rect 17083 14365 17092 14399
rect 17040 14356 17092 14365
rect 17868 14356 17920 14408
rect 18052 14399 18104 14408
rect 18052 14365 18061 14399
rect 18061 14365 18095 14399
rect 18095 14365 18104 14399
rect 18052 14356 18104 14365
rect 18512 14356 18564 14408
rect 19248 14399 19300 14408
rect 19248 14365 19257 14399
rect 19257 14365 19291 14399
rect 19291 14365 19300 14399
rect 19248 14356 19300 14365
rect 20168 14399 20220 14408
rect 20168 14365 20177 14399
rect 20177 14365 20211 14399
rect 20211 14365 20220 14399
rect 20168 14356 20220 14365
rect 21180 14399 21232 14408
rect 21180 14365 21189 14399
rect 21189 14365 21223 14399
rect 21223 14365 21232 14399
rect 21180 14356 21232 14365
rect 21640 14356 21692 14408
rect 22008 14399 22060 14408
rect 22008 14365 22017 14399
rect 22017 14365 22051 14399
rect 22051 14365 22060 14399
rect 22008 14356 22060 14365
rect 22652 14399 22704 14408
rect 22652 14365 22661 14399
rect 22661 14365 22695 14399
rect 22695 14365 22704 14399
rect 22652 14356 22704 14365
rect 23848 14399 23900 14408
rect 19064 14288 19116 14340
rect 15752 14220 15804 14272
rect 18420 14220 18472 14272
rect 18880 14220 18932 14272
rect 20352 14263 20404 14272
rect 20352 14229 20361 14263
rect 20361 14229 20395 14263
rect 20395 14229 20404 14263
rect 20352 14220 20404 14229
rect 20536 14288 20588 14340
rect 20996 14288 21048 14340
rect 22376 14288 22428 14340
rect 23848 14365 23857 14399
rect 23857 14365 23891 14399
rect 23891 14365 23900 14399
rect 23848 14356 23900 14365
rect 23940 14356 23992 14408
rect 20720 14220 20772 14272
rect 23388 14263 23440 14272
rect 23388 14229 23397 14263
rect 23397 14229 23431 14263
rect 23431 14229 23440 14263
rect 23388 14220 23440 14229
rect 25872 14288 25924 14340
rect 24492 14220 24544 14272
rect 28080 14220 28132 14272
rect 10214 14118 10266 14170
rect 10278 14118 10330 14170
rect 10342 14118 10394 14170
rect 10406 14118 10458 14170
rect 10470 14118 10522 14170
rect 19478 14118 19530 14170
rect 19542 14118 19594 14170
rect 19606 14118 19658 14170
rect 19670 14118 19722 14170
rect 19734 14118 19786 14170
rect 6920 14059 6972 14068
rect 6920 14025 6929 14059
rect 6929 14025 6963 14059
rect 6963 14025 6972 14059
rect 6920 14016 6972 14025
rect 8116 14016 8168 14068
rect 6552 13948 6604 14000
rect 6276 13880 6328 13932
rect 7104 13923 7156 13932
rect 7104 13889 7113 13923
rect 7113 13889 7147 13923
rect 7147 13889 7156 13923
rect 7104 13880 7156 13889
rect 8024 13948 8076 14000
rect 8484 13923 8536 13932
rect 1400 13855 1452 13864
rect 1400 13821 1409 13855
rect 1409 13821 1443 13855
rect 1443 13821 1452 13855
rect 1400 13812 1452 13821
rect 4436 13812 4488 13864
rect 6736 13812 6788 13864
rect 7012 13676 7064 13728
rect 8116 13812 8168 13864
rect 8484 13889 8493 13923
rect 8493 13889 8527 13923
rect 8527 13889 8536 13923
rect 8484 13880 8536 13889
rect 8576 13923 8628 13932
rect 8576 13889 8585 13923
rect 8585 13889 8619 13923
rect 8619 13889 8628 13923
rect 8944 13923 8996 13932
rect 8576 13880 8628 13889
rect 8944 13889 8953 13923
rect 8953 13889 8987 13923
rect 8987 13889 8996 13923
rect 8944 13880 8996 13889
rect 10140 13948 10192 14000
rect 9588 13880 9640 13932
rect 11704 13923 11756 13932
rect 11704 13889 11713 13923
rect 11713 13889 11747 13923
rect 11747 13889 11756 13923
rect 11704 13880 11756 13889
rect 12164 13923 12216 13932
rect 12164 13889 12173 13923
rect 12173 13889 12207 13923
rect 12207 13889 12216 13923
rect 12164 13880 12216 13889
rect 13084 14016 13136 14068
rect 13176 14059 13228 14068
rect 13176 14025 13185 14059
rect 13185 14025 13219 14059
rect 13219 14025 13228 14059
rect 13176 14016 13228 14025
rect 12440 13991 12492 14000
rect 12440 13957 12449 13991
rect 12449 13957 12483 13991
rect 12483 13957 12492 13991
rect 12440 13948 12492 13957
rect 15200 14016 15252 14068
rect 15384 14016 15436 14068
rect 15844 13948 15896 14000
rect 19248 14016 19300 14068
rect 20352 14016 20404 14068
rect 12532 13923 12584 13932
rect 12532 13889 12541 13923
rect 12541 13889 12575 13923
rect 12575 13889 12584 13923
rect 12532 13880 12584 13889
rect 13360 13880 13412 13932
rect 13728 13923 13780 13932
rect 13728 13889 13737 13923
rect 13737 13889 13771 13923
rect 13771 13889 13780 13923
rect 13728 13880 13780 13889
rect 8300 13812 8352 13864
rect 8208 13719 8260 13728
rect 8208 13685 8217 13719
rect 8217 13685 8251 13719
rect 8251 13685 8260 13719
rect 8208 13676 8260 13685
rect 12440 13744 12492 13796
rect 13636 13744 13688 13796
rect 13912 13923 13964 13932
rect 13912 13889 13921 13923
rect 13921 13889 13955 13923
rect 13955 13889 13964 13923
rect 13912 13880 13964 13889
rect 14464 13880 14516 13932
rect 15660 13880 15712 13932
rect 17040 13880 17092 13932
rect 17776 13923 17828 13932
rect 17776 13889 17785 13923
rect 17785 13889 17819 13923
rect 17819 13889 17828 13923
rect 17776 13880 17828 13889
rect 8392 13719 8444 13728
rect 8392 13685 8401 13719
rect 8401 13685 8435 13719
rect 8435 13685 8444 13719
rect 8392 13676 8444 13685
rect 9128 13676 9180 13728
rect 9496 13676 9548 13728
rect 10232 13676 10284 13728
rect 11704 13676 11756 13728
rect 12808 13719 12860 13728
rect 12808 13685 12817 13719
rect 12817 13685 12851 13719
rect 12851 13685 12860 13719
rect 12808 13676 12860 13685
rect 13728 13676 13780 13728
rect 16672 13855 16724 13864
rect 16672 13821 16681 13855
rect 16681 13821 16715 13855
rect 16715 13821 16724 13855
rect 16672 13812 16724 13821
rect 18328 13948 18380 14000
rect 18420 13923 18472 13932
rect 18420 13889 18429 13923
rect 18429 13889 18463 13923
rect 18463 13889 18472 13923
rect 18420 13880 18472 13889
rect 18880 13948 18932 14000
rect 20536 13991 20588 14000
rect 20536 13957 20545 13991
rect 20545 13957 20579 13991
rect 20579 13957 20588 13991
rect 20536 13948 20588 13957
rect 23388 13948 23440 14000
rect 19984 13880 20036 13932
rect 20904 13923 20956 13932
rect 20904 13889 20913 13923
rect 20913 13889 20947 13923
rect 20947 13889 20956 13923
rect 20904 13880 20956 13889
rect 21180 13880 21232 13932
rect 23572 13880 23624 13932
rect 24492 13880 24544 13932
rect 24952 13923 25004 13932
rect 24952 13889 24961 13923
rect 24961 13889 24995 13923
rect 24995 13889 25004 13923
rect 24952 13880 25004 13889
rect 25872 14016 25924 14068
rect 26056 14059 26108 14068
rect 26056 14025 26065 14059
rect 26065 14025 26099 14059
rect 26099 14025 26108 14059
rect 26056 14016 26108 14025
rect 26424 14059 26476 14068
rect 26424 14025 26433 14059
rect 26433 14025 26467 14059
rect 26467 14025 26476 14059
rect 26424 14016 26476 14025
rect 28264 13923 28316 13932
rect 28264 13889 28273 13923
rect 28273 13889 28307 13923
rect 28307 13889 28316 13923
rect 28264 13880 28316 13889
rect 16028 13744 16080 13796
rect 16396 13744 16448 13796
rect 14188 13676 14240 13728
rect 14648 13676 14700 13728
rect 17960 13719 18012 13728
rect 17960 13685 17969 13719
rect 17969 13685 18003 13719
rect 18003 13685 18012 13719
rect 17960 13676 18012 13685
rect 18144 13719 18196 13728
rect 18144 13685 18153 13719
rect 18153 13685 18187 13719
rect 18187 13685 18196 13719
rect 18144 13676 18196 13685
rect 18604 13676 18656 13728
rect 23940 13812 23992 13864
rect 23388 13744 23440 13796
rect 24676 13812 24728 13864
rect 25044 13812 25096 13864
rect 21732 13676 21784 13728
rect 22560 13676 22612 13728
rect 23664 13719 23716 13728
rect 23664 13685 23673 13719
rect 23673 13685 23707 13719
rect 23707 13685 23716 13719
rect 23664 13676 23716 13685
rect 25412 13676 25464 13728
rect 5582 13574 5634 13626
rect 5646 13574 5698 13626
rect 5710 13574 5762 13626
rect 5774 13574 5826 13626
rect 5838 13574 5890 13626
rect 14846 13574 14898 13626
rect 14910 13574 14962 13626
rect 14974 13574 15026 13626
rect 15038 13574 15090 13626
rect 15102 13574 15154 13626
rect 24110 13574 24162 13626
rect 24174 13574 24226 13626
rect 24238 13574 24290 13626
rect 24302 13574 24354 13626
rect 24366 13574 24418 13626
rect 6276 13515 6328 13524
rect 6276 13481 6285 13515
rect 6285 13481 6319 13515
rect 6319 13481 6328 13515
rect 6276 13472 6328 13481
rect 6552 13515 6604 13524
rect 6552 13481 6561 13515
rect 6561 13481 6595 13515
rect 6595 13481 6604 13515
rect 6552 13472 6604 13481
rect 7104 13472 7156 13524
rect 7932 13472 7984 13524
rect 8116 13472 8168 13524
rect 9588 13515 9640 13524
rect 7656 13404 7708 13456
rect 8208 13404 8260 13456
rect 6828 13336 6880 13388
rect 8392 13336 8444 13388
rect 9588 13481 9597 13515
rect 9597 13481 9631 13515
rect 9631 13481 9640 13515
rect 9588 13472 9640 13481
rect 9496 13404 9548 13456
rect 12164 13472 12216 13524
rect 13912 13472 13964 13524
rect 14280 13472 14332 13524
rect 15200 13472 15252 13524
rect 15568 13472 15620 13524
rect 16764 13472 16816 13524
rect 6736 13311 6788 13320
rect 6736 13277 6745 13311
rect 6745 13277 6779 13311
rect 6779 13277 6788 13311
rect 6736 13268 6788 13277
rect 7380 13268 7432 13320
rect 9128 13311 9180 13320
rect 9128 13277 9137 13311
rect 9137 13277 9171 13311
rect 9171 13277 9180 13311
rect 9128 13268 9180 13277
rect 11704 13336 11756 13388
rect 8484 13200 8536 13252
rect 8760 13200 8812 13252
rect 12072 13268 12124 13320
rect 12624 13311 12676 13320
rect 12624 13277 12631 13311
rect 12631 13277 12676 13311
rect 12624 13268 12676 13277
rect 13820 13404 13872 13456
rect 14740 13404 14792 13456
rect 16672 13404 16724 13456
rect 16028 13336 16080 13388
rect 16120 13336 16172 13388
rect 16856 13336 16908 13388
rect 17960 13472 18012 13524
rect 20076 13472 20128 13524
rect 20536 13472 20588 13524
rect 22008 13472 22060 13524
rect 23848 13515 23900 13524
rect 23848 13481 23857 13515
rect 23857 13481 23891 13515
rect 23891 13481 23900 13515
rect 23848 13472 23900 13481
rect 24952 13472 25004 13524
rect 13360 13311 13412 13320
rect 13360 13277 13369 13311
rect 13369 13277 13403 13311
rect 13403 13277 13412 13311
rect 13360 13268 13412 13277
rect 13636 13268 13688 13320
rect 15568 13268 15620 13320
rect 15752 13311 15804 13320
rect 15752 13277 15761 13311
rect 15761 13277 15795 13311
rect 15795 13277 15804 13311
rect 15752 13268 15804 13277
rect 16396 13311 16448 13320
rect 16396 13277 16405 13311
rect 16405 13277 16439 13311
rect 16439 13277 16448 13311
rect 16396 13268 16448 13277
rect 16580 13268 16632 13320
rect 20904 13404 20956 13456
rect 18052 13336 18104 13388
rect 22284 13336 22336 13388
rect 23388 13336 23440 13388
rect 24952 13336 25004 13388
rect 17408 13311 17460 13320
rect 17408 13277 17417 13311
rect 17417 13277 17451 13311
rect 17451 13277 17460 13311
rect 17408 13268 17460 13277
rect 10232 13243 10284 13252
rect 10232 13209 10241 13243
rect 10241 13209 10275 13243
rect 10275 13209 10284 13243
rect 10232 13200 10284 13209
rect 14188 13200 14240 13252
rect 7472 13132 7524 13184
rect 8208 13175 8260 13184
rect 8208 13141 8217 13175
rect 8217 13141 8251 13175
rect 8251 13141 8260 13175
rect 8208 13132 8260 13141
rect 8852 13132 8904 13184
rect 8944 13132 8996 13184
rect 11152 13132 11204 13184
rect 12900 13132 12952 13184
rect 13176 13132 13228 13184
rect 17040 13200 17092 13252
rect 15936 13175 15988 13184
rect 15936 13141 15945 13175
rect 15945 13141 15979 13175
rect 15979 13141 15988 13175
rect 15936 13132 15988 13141
rect 17224 13132 17276 13184
rect 17592 13311 17644 13320
rect 17592 13277 17601 13311
rect 17601 13277 17635 13311
rect 17635 13277 17644 13311
rect 17592 13268 17644 13277
rect 18420 13268 18472 13320
rect 18604 13311 18656 13320
rect 18604 13277 18613 13311
rect 18613 13277 18647 13311
rect 18647 13277 18656 13311
rect 18604 13268 18656 13277
rect 19248 13311 19300 13320
rect 19248 13277 19257 13311
rect 19257 13277 19291 13311
rect 19291 13277 19300 13311
rect 19248 13268 19300 13277
rect 17960 13200 18012 13252
rect 19892 13268 19944 13320
rect 21180 13311 21232 13320
rect 21180 13277 21189 13311
rect 21189 13277 21223 13311
rect 21223 13277 21232 13311
rect 21180 13268 21232 13277
rect 21732 13268 21784 13320
rect 22468 13268 22520 13320
rect 23296 13268 23348 13320
rect 23664 13311 23716 13320
rect 20352 13243 20404 13252
rect 20352 13209 20361 13243
rect 20361 13209 20395 13243
rect 20395 13209 20404 13243
rect 20352 13200 20404 13209
rect 23664 13277 23673 13311
rect 23673 13277 23707 13311
rect 23707 13277 23716 13311
rect 23664 13268 23716 13277
rect 23940 13268 23992 13320
rect 24768 13268 24820 13320
rect 18328 13132 18380 13184
rect 20720 13175 20772 13184
rect 20720 13141 20729 13175
rect 20729 13141 20763 13175
rect 20763 13141 20772 13175
rect 20720 13132 20772 13141
rect 21180 13132 21232 13184
rect 21640 13132 21692 13184
rect 24676 13200 24728 13252
rect 22652 13175 22704 13184
rect 22652 13141 22661 13175
rect 22661 13141 22695 13175
rect 22695 13141 22704 13175
rect 22652 13132 22704 13141
rect 24860 13175 24912 13184
rect 24860 13141 24869 13175
rect 24869 13141 24903 13175
rect 24903 13141 24912 13175
rect 24860 13132 24912 13141
rect 25320 13132 25372 13184
rect 25596 13200 25648 13252
rect 25872 13132 25924 13184
rect 10214 13030 10266 13082
rect 10278 13030 10330 13082
rect 10342 13030 10394 13082
rect 10406 13030 10458 13082
rect 10470 13030 10522 13082
rect 19478 13030 19530 13082
rect 19542 13030 19594 13082
rect 19606 13030 19658 13082
rect 19670 13030 19722 13082
rect 19734 13030 19786 13082
rect 6736 12928 6788 12980
rect 7472 12971 7524 12980
rect 7104 12860 7156 12912
rect 7472 12937 7481 12971
rect 7481 12937 7515 12971
rect 7515 12937 7524 12971
rect 7472 12928 7524 12937
rect 7932 12971 7984 12980
rect 7932 12937 7941 12971
rect 7941 12937 7975 12971
rect 7975 12937 7984 12971
rect 7932 12928 7984 12937
rect 8760 12928 8812 12980
rect 9496 12928 9548 12980
rect 12532 12928 12584 12980
rect 13636 12928 13688 12980
rect 15660 12971 15712 12980
rect 15660 12937 15669 12971
rect 15669 12937 15703 12971
rect 15703 12937 15712 12971
rect 15660 12928 15712 12937
rect 16948 12928 17000 12980
rect 17408 12928 17460 12980
rect 18972 12928 19024 12980
rect 19248 12928 19300 12980
rect 20444 12928 20496 12980
rect 22744 12928 22796 12980
rect 24032 12971 24084 12980
rect 24032 12937 24041 12971
rect 24041 12937 24075 12971
rect 24075 12937 24084 12971
rect 24032 12928 24084 12937
rect 25596 12971 25648 12980
rect 25596 12937 25605 12971
rect 25605 12937 25639 12971
rect 25639 12937 25648 12971
rect 25596 12928 25648 12937
rect 8944 12903 8996 12912
rect 4436 12835 4488 12844
rect 4436 12801 4445 12835
rect 4445 12801 4479 12835
rect 4479 12801 4488 12835
rect 4436 12792 4488 12801
rect 5908 12792 5960 12844
rect 7472 12835 7524 12844
rect 7472 12801 7481 12835
rect 7481 12801 7515 12835
rect 7515 12801 7524 12835
rect 7472 12792 7524 12801
rect 8944 12869 8955 12903
rect 8955 12869 8996 12903
rect 8944 12860 8996 12869
rect 8484 12792 8536 12844
rect 12348 12860 12400 12912
rect 14372 12903 14424 12912
rect 14372 12869 14381 12903
rect 14381 12869 14415 12903
rect 14415 12869 14424 12903
rect 14372 12860 14424 12869
rect 8024 12724 8076 12776
rect 8668 12724 8720 12776
rect 9680 12767 9732 12776
rect 6092 12588 6144 12640
rect 6828 12631 6880 12640
rect 6828 12597 6837 12631
rect 6837 12597 6871 12631
rect 6871 12597 6880 12631
rect 6828 12588 6880 12597
rect 7012 12631 7064 12640
rect 7012 12597 7021 12631
rect 7021 12597 7055 12631
rect 7055 12597 7064 12631
rect 7012 12588 7064 12597
rect 8208 12588 8260 12640
rect 9680 12733 9689 12767
rect 9689 12733 9723 12767
rect 9723 12733 9732 12767
rect 9680 12724 9732 12733
rect 9864 12724 9916 12776
rect 13176 12792 13228 12844
rect 14188 12792 14240 12844
rect 15936 12860 15988 12912
rect 16396 12860 16448 12912
rect 11612 12767 11664 12776
rect 11612 12733 11621 12767
rect 11621 12733 11655 12767
rect 11655 12733 11664 12767
rect 11612 12724 11664 12733
rect 12072 12767 12124 12776
rect 12072 12733 12081 12767
rect 12081 12733 12115 12767
rect 12115 12733 12124 12767
rect 12072 12724 12124 12733
rect 14464 12724 14516 12776
rect 14648 12724 14700 12776
rect 15292 12792 15344 12844
rect 15844 12792 15896 12844
rect 16672 12792 16724 12844
rect 15568 12724 15620 12776
rect 13360 12656 13412 12708
rect 14096 12656 14148 12708
rect 16672 12656 16724 12708
rect 17500 12792 17552 12844
rect 20904 12860 20956 12912
rect 24584 12860 24636 12912
rect 16856 12724 16908 12776
rect 18880 12724 18932 12776
rect 19340 12724 19392 12776
rect 10968 12631 11020 12640
rect 10968 12597 10977 12631
rect 10977 12597 11011 12631
rect 11011 12597 11020 12631
rect 10968 12588 11020 12597
rect 12716 12588 12768 12640
rect 14648 12588 14700 12640
rect 16120 12588 16172 12640
rect 16580 12588 16632 12640
rect 17224 12588 17276 12640
rect 17316 12588 17368 12640
rect 18880 12631 18932 12640
rect 18880 12597 18889 12631
rect 18889 12597 18923 12631
rect 18923 12597 18932 12631
rect 18880 12588 18932 12597
rect 19340 12588 19392 12640
rect 20168 12792 20220 12844
rect 21088 12792 21140 12844
rect 21180 12792 21232 12844
rect 23020 12792 23072 12844
rect 25412 12835 25464 12844
rect 25412 12801 25421 12835
rect 25421 12801 25455 12835
rect 25455 12801 25464 12835
rect 25412 12792 25464 12801
rect 26056 12835 26108 12844
rect 26056 12801 26065 12835
rect 26065 12801 26099 12835
rect 26099 12801 26108 12835
rect 26056 12792 26108 12801
rect 20076 12767 20128 12776
rect 20076 12733 20085 12767
rect 20085 12733 20119 12767
rect 20119 12733 20128 12767
rect 20076 12724 20128 12733
rect 24860 12767 24912 12776
rect 22284 12656 22336 12708
rect 21456 12631 21508 12640
rect 21456 12597 21465 12631
rect 21465 12597 21499 12631
rect 21499 12597 21508 12631
rect 21456 12588 21508 12597
rect 24860 12733 24869 12767
rect 24869 12733 24903 12767
rect 24903 12733 24912 12767
rect 24860 12724 24912 12733
rect 24952 12767 25004 12776
rect 24952 12733 24961 12767
rect 24961 12733 24995 12767
rect 24995 12733 25004 12767
rect 24952 12724 25004 12733
rect 23480 12588 23532 12640
rect 23756 12631 23808 12640
rect 23756 12597 23765 12631
rect 23765 12597 23799 12631
rect 23799 12597 23808 12631
rect 23756 12588 23808 12597
rect 24584 12588 24636 12640
rect 25688 12588 25740 12640
rect 28356 12631 28408 12640
rect 28356 12597 28365 12631
rect 28365 12597 28399 12631
rect 28399 12597 28408 12631
rect 28356 12588 28408 12597
rect 5582 12486 5634 12538
rect 5646 12486 5698 12538
rect 5710 12486 5762 12538
rect 5774 12486 5826 12538
rect 5838 12486 5890 12538
rect 14846 12486 14898 12538
rect 14910 12486 14962 12538
rect 14974 12486 15026 12538
rect 15038 12486 15090 12538
rect 15102 12486 15154 12538
rect 24110 12486 24162 12538
rect 24174 12486 24226 12538
rect 24238 12486 24290 12538
rect 24302 12486 24354 12538
rect 24366 12486 24418 12538
rect 5908 12384 5960 12436
rect 6920 12384 6972 12436
rect 7012 12384 7064 12436
rect 8392 12384 8444 12436
rect 8576 12427 8628 12436
rect 8576 12393 8585 12427
rect 8585 12393 8619 12427
rect 8619 12393 8628 12427
rect 8576 12384 8628 12393
rect 9680 12384 9732 12436
rect 10600 12427 10652 12436
rect 6644 12316 6696 12368
rect 7380 12316 7432 12368
rect 8024 12316 8076 12368
rect 8116 12316 8168 12368
rect 6828 12248 6880 12300
rect 6000 12223 6052 12232
rect 6000 12189 6009 12223
rect 6009 12189 6043 12223
rect 6043 12189 6052 12223
rect 6000 12180 6052 12189
rect 6644 12180 6696 12232
rect 7564 12180 7616 12232
rect 9864 12316 9916 12368
rect 10048 12316 10100 12368
rect 10600 12393 10609 12427
rect 10609 12393 10643 12427
rect 10643 12393 10652 12427
rect 10600 12384 10652 12393
rect 11612 12384 11664 12436
rect 12348 12427 12400 12436
rect 12348 12393 12357 12427
rect 12357 12393 12391 12427
rect 12391 12393 12400 12427
rect 12348 12384 12400 12393
rect 15384 12384 15436 12436
rect 16580 12384 16632 12436
rect 20352 12384 20404 12436
rect 21824 12384 21876 12436
rect 23940 12384 23992 12436
rect 26056 12384 26108 12436
rect 8852 12248 8904 12300
rect 14556 12316 14608 12368
rect 14832 12316 14884 12368
rect 9680 12180 9732 12232
rect 11980 12291 12032 12300
rect 11980 12257 11989 12291
rect 11989 12257 12023 12291
rect 12023 12257 12032 12291
rect 11980 12248 12032 12257
rect 11152 12180 11204 12232
rect 13636 12180 13688 12232
rect 13820 12180 13872 12232
rect 15200 12248 15252 12300
rect 14648 12223 14700 12232
rect 14648 12189 14657 12223
rect 14657 12189 14691 12223
rect 14691 12189 14700 12223
rect 14648 12180 14700 12189
rect 14832 12223 14884 12232
rect 14832 12189 14841 12223
rect 14841 12189 14875 12223
rect 14875 12189 14884 12223
rect 14832 12180 14884 12189
rect 6092 12112 6144 12164
rect 6552 12155 6604 12164
rect 6552 12121 6561 12155
rect 6561 12121 6595 12155
rect 6595 12121 6604 12155
rect 6552 12112 6604 12121
rect 6736 12155 6788 12164
rect 6736 12121 6761 12155
rect 6761 12121 6788 12155
rect 7472 12155 7524 12164
rect 6736 12112 6788 12121
rect 7472 12121 7481 12155
rect 7481 12121 7515 12155
rect 7515 12121 7524 12155
rect 7472 12112 7524 12121
rect 8208 12112 8260 12164
rect 7012 12044 7064 12096
rect 7748 12044 7800 12096
rect 8024 12044 8076 12096
rect 9312 12155 9364 12164
rect 9312 12121 9321 12155
rect 9321 12121 9355 12155
rect 9355 12121 9364 12155
rect 9312 12112 9364 12121
rect 10876 12112 10928 12164
rect 15568 12223 15620 12232
rect 15568 12189 15577 12223
rect 15577 12189 15611 12223
rect 15611 12189 15620 12223
rect 17592 12316 17644 12368
rect 15568 12180 15620 12189
rect 16120 12223 16172 12232
rect 16120 12189 16129 12223
rect 16129 12189 16163 12223
rect 16163 12189 16172 12223
rect 17040 12248 17092 12300
rect 17224 12248 17276 12300
rect 16120 12180 16172 12189
rect 16396 12223 16448 12232
rect 16396 12189 16405 12223
rect 16405 12189 16439 12223
rect 16439 12189 16448 12223
rect 16396 12180 16448 12189
rect 17316 12223 17368 12232
rect 17316 12189 17325 12223
rect 17325 12189 17359 12223
rect 17359 12189 17368 12223
rect 17316 12180 17368 12189
rect 21180 12248 21232 12300
rect 17500 12223 17552 12232
rect 17500 12189 17509 12223
rect 17509 12189 17543 12223
rect 17543 12189 17552 12223
rect 17500 12180 17552 12189
rect 19984 12180 20036 12232
rect 20812 12223 20864 12232
rect 20812 12189 20821 12223
rect 20821 12189 20855 12223
rect 20855 12189 20864 12223
rect 20812 12180 20864 12189
rect 21364 12180 21416 12232
rect 22192 12248 22244 12300
rect 22284 12248 22336 12300
rect 25044 12316 25096 12368
rect 21640 12223 21692 12232
rect 21640 12189 21649 12223
rect 21649 12189 21683 12223
rect 21683 12189 21692 12223
rect 21640 12180 21692 12189
rect 24676 12248 24728 12300
rect 18052 12112 18104 12164
rect 19892 12155 19944 12164
rect 19892 12121 19901 12155
rect 19901 12121 19935 12155
rect 19935 12121 19944 12155
rect 19892 12112 19944 12121
rect 8668 12044 8720 12096
rect 14188 12087 14240 12096
rect 14188 12053 14197 12087
rect 14197 12053 14231 12087
rect 14231 12053 14240 12087
rect 14188 12044 14240 12053
rect 16580 12087 16632 12096
rect 16580 12053 16589 12087
rect 16589 12053 16623 12087
rect 16623 12053 16632 12087
rect 16580 12044 16632 12053
rect 17776 12087 17828 12096
rect 17776 12053 17785 12087
rect 17785 12053 17819 12087
rect 17819 12053 17828 12087
rect 17776 12044 17828 12053
rect 19340 12087 19392 12096
rect 19340 12053 19349 12087
rect 19349 12053 19383 12087
rect 19383 12053 19392 12087
rect 19340 12044 19392 12053
rect 21456 12044 21508 12096
rect 21916 12087 21968 12096
rect 21916 12053 21925 12087
rect 21925 12053 21959 12087
rect 21959 12053 21968 12087
rect 21916 12044 21968 12053
rect 23572 12180 23624 12232
rect 23756 12180 23808 12232
rect 24032 12223 24084 12232
rect 24032 12189 24041 12223
rect 24041 12189 24075 12223
rect 24075 12189 24084 12223
rect 24032 12180 24084 12189
rect 24584 12223 24636 12232
rect 24584 12189 24593 12223
rect 24593 12189 24627 12223
rect 24627 12189 24636 12223
rect 24584 12180 24636 12189
rect 24768 12180 24820 12232
rect 22560 12155 22612 12164
rect 22560 12121 22569 12155
rect 22569 12121 22603 12155
rect 22603 12121 22612 12155
rect 22560 12112 22612 12121
rect 23572 12044 23624 12096
rect 23848 12087 23900 12096
rect 23848 12053 23857 12087
rect 23857 12053 23891 12087
rect 23891 12053 23900 12087
rect 23848 12044 23900 12053
rect 25688 12155 25740 12164
rect 25688 12121 25722 12155
rect 25722 12121 25740 12155
rect 25688 12112 25740 12121
rect 25780 12044 25832 12096
rect 25964 12044 26016 12096
rect 10214 11942 10266 11994
rect 10278 11942 10330 11994
rect 10342 11942 10394 11994
rect 10406 11942 10458 11994
rect 10470 11942 10522 11994
rect 19478 11942 19530 11994
rect 19542 11942 19594 11994
rect 19606 11942 19658 11994
rect 19670 11942 19722 11994
rect 19734 11942 19786 11994
rect 4528 11704 4580 11756
rect 7104 11840 7156 11892
rect 7840 11840 7892 11892
rect 10692 11840 10744 11892
rect 10876 11883 10928 11892
rect 10876 11849 10885 11883
rect 10885 11849 10919 11883
rect 10919 11849 10928 11883
rect 10876 11840 10928 11849
rect 11152 11840 11204 11892
rect 12256 11840 12308 11892
rect 12992 11883 13044 11892
rect 12992 11849 13001 11883
rect 13001 11849 13035 11883
rect 13035 11849 13044 11883
rect 12992 11840 13044 11849
rect 15844 11883 15896 11892
rect 15844 11849 15853 11883
rect 15853 11849 15887 11883
rect 15887 11849 15896 11883
rect 15844 11840 15896 11849
rect 17868 11840 17920 11892
rect 20444 11883 20496 11892
rect 6000 11704 6052 11756
rect 7472 11772 7524 11824
rect 14188 11772 14240 11824
rect 7012 11636 7064 11688
rect 7380 11704 7432 11756
rect 7656 11704 7708 11756
rect 8392 11704 8444 11756
rect 7564 11636 7616 11688
rect 8208 11636 8260 11688
rect 8760 11636 8812 11688
rect 7656 11568 7708 11620
rect 9680 11704 9732 11756
rect 10048 11704 10100 11756
rect 10232 11747 10284 11756
rect 10232 11713 10241 11747
rect 10241 11713 10275 11747
rect 10275 11713 10284 11747
rect 10232 11704 10284 11713
rect 10324 11704 10376 11756
rect 10324 11568 10376 11620
rect 5448 11500 5500 11552
rect 6828 11500 6880 11552
rect 9772 11543 9824 11552
rect 9772 11509 9781 11543
rect 9781 11509 9815 11543
rect 9815 11509 9824 11543
rect 9772 11500 9824 11509
rect 10140 11500 10192 11552
rect 10600 11747 10652 11756
rect 10600 11713 10609 11747
rect 10609 11713 10643 11747
rect 10643 11713 10652 11747
rect 12072 11747 12124 11756
rect 10600 11704 10652 11713
rect 12072 11713 12081 11747
rect 12081 11713 12115 11747
rect 12115 11713 12124 11747
rect 12072 11704 12124 11713
rect 12256 11704 12308 11756
rect 13636 11704 13688 11756
rect 16580 11772 16632 11824
rect 20444 11849 20453 11883
rect 20453 11849 20487 11883
rect 20487 11849 20496 11883
rect 20444 11840 20496 11849
rect 20904 11840 20956 11892
rect 21088 11883 21140 11892
rect 21088 11849 21097 11883
rect 21097 11849 21131 11883
rect 21131 11849 21140 11883
rect 21088 11840 21140 11849
rect 23020 11883 23072 11892
rect 13728 11636 13780 11688
rect 15292 11704 15344 11756
rect 10600 11500 10652 11552
rect 13176 11568 13228 11620
rect 17040 11704 17092 11756
rect 20996 11772 21048 11824
rect 21916 11772 21968 11824
rect 18052 11679 18104 11688
rect 18052 11645 18061 11679
rect 18061 11645 18095 11679
rect 18095 11645 18104 11679
rect 18052 11636 18104 11645
rect 19984 11704 20036 11756
rect 20720 11704 20772 11756
rect 22100 11747 22152 11756
rect 22100 11713 22109 11747
rect 22109 11713 22143 11747
rect 22143 11713 22152 11747
rect 22100 11704 22152 11713
rect 22376 11704 22428 11756
rect 23020 11849 23029 11883
rect 23029 11849 23063 11883
rect 23063 11849 23072 11883
rect 23020 11840 23072 11849
rect 24492 11883 24544 11892
rect 24492 11849 24501 11883
rect 24501 11849 24535 11883
rect 24535 11849 24544 11883
rect 24492 11840 24544 11849
rect 24860 11840 24912 11892
rect 25964 11883 26016 11892
rect 25964 11849 25973 11883
rect 25973 11849 26007 11883
rect 26007 11849 26016 11883
rect 25964 11840 26016 11849
rect 20260 11636 20312 11688
rect 20536 11568 20588 11620
rect 21180 11636 21232 11688
rect 11980 11500 12032 11552
rect 13268 11500 13320 11552
rect 13820 11543 13872 11552
rect 13820 11509 13829 11543
rect 13829 11509 13863 11543
rect 13863 11509 13872 11543
rect 13820 11500 13872 11509
rect 13912 11500 13964 11552
rect 16120 11500 16172 11552
rect 18512 11500 18564 11552
rect 18972 11543 19024 11552
rect 18972 11509 18981 11543
rect 18981 11509 19015 11543
rect 19015 11509 19024 11543
rect 18972 11500 19024 11509
rect 19156 11500 19208 11552
rect 20352 11500 20404 11552
rect 21180 11500 21232 11552
rect 23480 11704 23532 11756
rect 24768 11772 24820 11824
rect 25320 11772 25372 11824
rect 25136 11704 25188 11756
rect 25504 11636 25556 11688
rect 26056 11679 26108 11688
rect 26056 11645 26065 11679
rect 26065 11645 26099 11679
rect 26099 11645 26108 11679
rect 26056 11636 26108 11645
rect 28264 11747 28316 11756
rect 28264 11713 28273 11747
rect 28273 11713 28307 11747
rect 28307 11713 28316 11747
rect 28264 11704 28316 11713
rect 22560 11543 22612 11552
rect 22560 11509 22569 11543
rect 22569 11509 22603 11543
rect 22603 11509 22612 11543
rect 22560 11500 22612 11509
rect 23572 11500 23624 11552
rect 25044 11500 25096 11552
rect 5582 11398 5634 11450
rect 5646 11398 5698 11450
rect 5710 11398 5762 11450
rect 5774 11398 5826 11450
rect 5838 11398 5890 11450
rect 14846 11398 14898 11450
rect 14910 11398 14962 11450
rect 14974 11398 15026 11450
rect 15038 11398 15090 11450
rect 15102 11398 15154 11450
rect 24110 11398 24162 11450
rect 24174 11398 24226 11450
rect 24238 11398 24290 11450
rect 24302 11398 24354 11450
rect 24366 11398 24418 11450
rect 4528 11339 4580 11348
rect 4528 11305 4537 11339
rect 4537 11305 4571 11339
rect 4571 11305 4580 11339
rect 4528 11296 4580 11305
rect 6552 11296 6604 11348
rect 7012 11296 7064 11348
rect 7656 11271 7708 11280
rect 7196 11160 7248 11212
rect 7656 11237 7665 11271
rect 7665 11237 7699 11271
rect 7699 11237 7708 11271
rect 7656 11228 7708 11237
rect 9312 11296 9364 11348
rect 9772 11296 9824 11348
rect 10416 11296 10468 11348
rect 12808 11296 12860 11348
rect 15476 11296 15528 11348
rect 15660 11296 15712 11348
rect 17040 11339 17092 11348
rect 17040 11305 17049 11339
rect 17049 11305 17083 11339
rect 17083 11305 17092 11339
rect 17040 11296 17092 11305
rect 17500 11296 17552 11348
rect 20812 11296 20864 11348
rect 20996 11339 21048 11348
rect 20996 11305 21005 11339
rect 21005 11305 21039 11339
rect 21039 11305 21048 11339
rect 20996 11296 21048 11305
rect 22100 11296 22152 11348
rect 26516 11296 26568 11348
rect 10692 11228 10744 11280
rect 5908 11135 5960 11144
rect 5908 11101 5917 11135
rect 5917 11101 5951 11135
rect 5951 11101 5960 11135
rect 5908 11092 5960 11101
rect 5540 11024 5592 11076
rect 6828 11067 6880 11076
rect 6828 11033 6837 11067
rect 6837 11033 6871 11067
rect 6871 11033 6880 11067
rect 6828 11024 6880 11033
rect 7104 11135 7156 11144
rect 7104 11101 7113 11135
rect 7113 11101 7147 11135
rect 7147 11101 7156 11135
rect 7104 11092 7156 11101
rect 7748 11135 7800 11144
rect 7748 11101 7757 11135
rect 7757 11101 7791 11135
rect 7791 11101 7800 11135
rect 7748 11092 7800 11101
rect 8116 11135 8168 11144
rect 8116 11101 8125 11135
rect 8125 11101 8159 11135
rect 8159 11101 8168 11135
rect 8116 11092 8168 11101
rect 8208 11135 8260 11144
rect 8208 11101 8217 11135
rect 8217 11101 8251 11135
rect 8251 11101 8260 11135
rect 8208 11092 8260 11101
rect 8852 11092 8904 11144
rect 8300 11024 8352 11076
rect 8944 11067 8996 11076
rect 8944 11033 8953 11067
rect 8953 11033 8987 11067
rect 8987 11033 8996 11067
rect 8944 11024 8996 11033
rect 12072 11160 12124 11212
rect 9496 11135 9548 11144
rect 9496 11101 9505 11135
rect 9505 11101 9539 11135
rect 9539 11101 9548 11135
rect 9496 11092 9548 11101
rect 9864 11092 9916 11144
rect 10600 11135 10652 11144
rect 10600 11101 10609 11135
rect 10609 11101 10643 11135
rect 10643 11101 10652 11135
rect 10600 11092 10652 11101
rect 10784 11135 10836 11144
rect 10784 11101 10793 11135
rect 10793 11101 10827 11135
rect 10827 11101 10836 11135
rect 10784 11092 10836 11101
rect 10140 11024 10192 11076
rect 10784 10956 10836 11008
rect 10968 11135 11020 11144
rect 10968 11101 10977 11135
rect 10977 11101 11011 11135
rect 11011 11101 11020 11135
rect 14372 11271 14424 11280
rect 14372 11237 14381 11271
rect 14381 11237 14415 11271
rect 14415 11237 14424 11271
rect 14372 11228 14424 11237
rect 14556 11228 14608 11280
rect 16304 11228 16356 11280
rect 16856 11228 16908 11280
rect 24032 11228 24084 11280
rect 15016 11203 15068 11212
rect 15016 11169 15025 11203
rect 15025 11169 15059 11203
rect 15059 11169 15068 11203
rect 15016 11160 15068 11169
rect 15200 11160 15252 11212
rect 15660 11160 15712 11212
rect 10968 11092 11020 11101
rect 12900 11092 12952 11144
rect 13084 11135 13136 11144
rect 13084 11101 13093 11135
rect 13093 11101 13127 11135
rect 13127 11101 13136 11135
rect 13084 11092 13136 11101
rect 13268 11135 13320 11144
rect 13268 11101 13277 11135
rect 13277 11101 13311 11135
rect 13311 11101 13320 11135
rect 13268 11092 13320 11101
rect 13452 11135 13504 11144
rect 13452 11101 13461 11135
rect 13461 11101 13495 11135
rect 13495 11101 13504 11135
rect 13452 11092 13504 11101
rect 14280 11092 14332 11144
rect 14648 11092 14700 11144
rect 11152 11024 11204 11076
rect 12992 11024 13044 11076
rect 13360 11067 13412 11076
rect 13360 11033 13369 11067
rect 13369 11033 13403 11067
rect 13403 11033 13412 11067
rect 13360 11024 13412 11033
rect 13912 11024 13964 11076
rect 15200 11067 15252 11076
rect 15200 11033 15209 11067
rect 15209 11033 15243 11067
rect 15243 11033 15252 11067
rect 15200 11024 15252 11033
rect 16120 11067 16172 11076
rect 16120 11033 16129 11067
rect 16129 11033 16163 11067
rect 16163 11033 16172 11067
rect 16120 11024 16172 11033
rect 11244 10999 11296 11008
rect 11244 10965 11253 10999
rect 11253 10965 11287 10999
rect 11287 10965 11296 10999
rect 11244 10956 11296 10965
rect 12072 10999 12124 11008
rect 12072 10965 12081 10999
rect 12081 10965 12115 10999
rect 12115 10965 12124 10999
rect 12072 10956 12124 10965
rect 18052 11092 18104 11144
rect 19248 11092 19300 11144
rect 23572 11160 23624 11212
rect 25044 11203 25096 11212
rect 25044 11169 25053 11203
rect 25053 11169 25087 11203
rect 25087 11169 25096 11203
rect 25044 11160 25096 11169
rect 24952 11092 25004 11144
rect 25136 11135 25188 11144
rect 25136 11101 25145 11135
rect 25145 11101 25179 11135
rect 25179 11101 25188 11135
rect 25136 11092 25188 11101
rect 25780 11135 25832 11144
rect 25780 11101 25789 11135
rect 25789 11101 25823 11135
rect 25823 11101 25832 11135
rect 25780 11092 25832 11101
rect 26332 11092 26384 11144
rect 17776 11024 17828 11076
rect 18972 11024 19024 11076
rect 20076 11024 20128 11076
rect 22560 11024 22612 11076
rect 22468 10956 22520 11008
rect 26424 11024 26476 11076
rect 10214 10854 10266 10906
rect 10278 10854 10330 10906
rect 10342 10854 10394 10906
rect 10406 10854 10458 10906
rect 10470 10854 10522 10906
rect 19478 10854 19530 10906
rect 19542 10854 19594 10906
rect 19606 10854 19658 10906
rect 19670 10854 19722 10906
rect 19734 10854 19786 10906
rect 7840 10795 7892 10804
rect 7840 10761 7849 10795
rect 7849 10761 7883 10795
rect 7883 10761 7892 10795
rect 7840 10752 7892 10761
rect 8116 10752 8168 10804
rect 10876 10795 10928 10804
rect 6000 10616 6052 10668
rect 7196 10684 7248 10736
rect 10876 10761 10885 10795
rect 10885 10761 10919 10795
rect 10919 10761 10928 10795
rect 10876 10752 10928 10761
rect 10968 10752 11020 10804
rect 9680 10684 9732 10736
rect 7104 10659 7156 10668
rect 7104 10625 7113 10659
rect 7113 10625 7147 10659
rect 7147 10625 7156 10659
rect 7104 10616 7156 10625
rect 7472 10616 7524 10668
rect 7748 10659 7800 10668
rect 7748 10625 7757 10659
rect 7757 10625 7791 10659
rect 7791 10625 7800 10659
rect 7748 10616 7800 10625
rect 8668 10659 8720 10668
rect 8668 10625 8677 10659
rect 8677 10625 8711 10659
rect 8711 10625 8720 10659
rect 8668 10616 8720 10625
rect 8944 10616 8996 10668
rect 10140 10616 10192 10668
rect 11244 10684 11296 10736
rect 11980 10684 12032 10736
rect 14188 10752 14240 10804
rect 16672 10752 16724 10804
rect 14372 10684 14424 10736
rect 19248 10795 19300 10804
rect 19248 10761 19257 10795
rect 19257 10761 19291 10795
rect 19291 10761 19300 10795
rect 19248 10752 19300 10761
rect 20260 10752 20312 10804
rect 20996 10752 21048 10804
rect 26424 10795 26476 10804
rect 26424 10761 26433 10795
rect 26433 10761 26467 10795
rect 26467 10761 26476 10795
rect 26424 10752 26476 10761
rect 18328 10684 18380 10736
rect 13268 10616 13320 10668
rect 15292 10659 15344 10668
rect 15292 10625 15301 10659
rect 15301 10625 15335 10659
rect 15335 10625 15344 10659
rect 15292 10616 15344 10625
rect 21180 10684 21232 10736
rect 21364 10727 21416 10736
rect 21364 10693 21373 10727
rect 21373 10693 21407 10727
rect 21407 10693 21416 10727
rect 21364 10684 21416 10693
rect 22468 10727 22520 10736
rect 22468 10693 22477 10727
rect 22477 10693 22511 10727
rect 22511 10693 22520 10727
rect 22468 10684 22520 10693
rect 23848 10684 23900 10736
rect 19892 10659 19944 10668
rect 19892 10625 19901 10659
rect 19901 10625 19935 10659
rect 19935 10625 19944 10659
rect 19892 10616 19944 10625
rect 20076 10659 20128 10668
rect 20076 10625 20085 10659
rect 20085 10625 20119 10659
rect 20119 10625 20128 10659
rect 20076 10616 20128 10625
rect 20352 10659 20404 10668
rect 20352 10625 20361 10659
rect 20361 10625 20395 10659
rect 20395 10625 20404 10659
rect 20352 10616 20404 10625
rect 6920 10480 6972 10532
rect 12808 10480 12860 10532
rect 13912 10548 13964 10600
rect 20904 10616 20956 10668
rect 21456 10616 21508 10668
rect 23480 10659 23532 10668
rect 22560 10591 22612 10600
rect 13544 10480 13596 10532
rect 1400 10455 1452 10464
rect 1400 10421 1409 10455
rect 1409 10421 1443 10455
rect 1443 10421 1452 10455
rect 1400 10412 1452 10421
rect 5448 10455 5500 10464
rect 5448 10421 5457 10455
rect 5457 10421 5491 10455
rect 5491 10421 5500 10455
rect 5448 10412 5500 10421
rect 6828 10455 6880 10464
rect 6828 10421 6837 10455
rect 6837 10421 6871 10455
rect 6871 10421 6880 10455
rect 6828 10412 6880 10421
rect 7104 10412 7156 10464
rect 7564 10412 7616 10464
rect 9036 10412 9088 10464
rect 11152 10412 11204 10464
rect 14096 10412 14148 10464
rect 14464 10412 14516 10464
rect 15200 10412 15252 10464
rect 15844 10412 15896 10464
rect 22560 10557 22569 10591
rect 22569 10557 22603 10591
rect 22603 10557 22612 10591
rect 22560 10548 22612 10557
rect 19432 10480 19484 10532
rect 20352 10480 20404 10532
rect 19340 10412 19392 10464
rect 21916 10412 21968 10464
rect 23020 10455 23072 10464
rect 23020 10421 23029 10455
rect 23029 10421 23063 10455
rect 23063 10421 23072 10455
rect 23020 10412 23072 10421
rect 23480 10625 23489 10659
rect 23489 10625 23523 10659
rect 23523 10625 23532 10659
rect 23480 10616 23532 10625
rect 26516 10616 26568 10668
rect 28080 10659 28132 10668
rect 28080 10625 28089 10659
rect 28089 10625 28123 10659
rect 28123 10625 28132 10659
rect 28080 10616 28132 10625
rect 25504 10591 25556 10600
rect 25504 10557 25513 10591
rect 25513 10557 25547 10591
rect 25547 10557 25556 10591
rect 25504 10548 25556 10557
rect 25688 10591 25740 10600
rect 25688 10557 25697 10591
rect 25697 10557 25731 10591
rect 25731 10557 25740 10591
rect 25688 10548 25740 10557
rect 25136 10480 25188 10532
rect 24676 10412 24728 10464
rect 26148 10455 26200 10464
rect 26148 10421 26157 10455
rect 26157 10421 26191 10455
rect 26191 10421 26200 10455
rect 26148 10412 26200 10421
rect 28264 10455 28316 10464
rect 28264 10421 28273 10455
rect 28273 10421 28307 10455
rect 28307 10421 28316 10455
rect 28264 10412 28316 10421
rect 5582 10310 5634 10362
rect 5646 10310 5698 10362
rect 5710 10310 5762 10362
rect 5774 10310 5826 10362
rect 5838 10310 5890 10362
rect 14846 10310 14898 10362
rect 14910 10310 14962 10362
rect 14974 10310 15026 10362
rect 15038 10310 15090 10362
rect 15102 10310 15154 10362
rect 24110 10310 24162 10362
rect 24174 10310 24226 10362
rect 24238 10310 24290 10362
rect 24302 10310 24354 10362
rect 24366 10310 24418 10362
rect 7288 10251 7340 10260
rect 7288 10217 7297 10251
rect 7297 10217 7331 10251
rect 7331 10217 7340 10251
rect 7288 10208 7340 10217
rect 8392 10208 8444 10260
rect 9036 10208 9088 10260
rect 6828 10140 6880 10192
rect 7748 10072 7800 10124
rect 9128 10115 9180 10124
rect 9128 10081 9137 10115
rect 9137 10081 9171 10115
rect 9171 10081 9180 10115
rect 9128 10072 9180 10081
rect 10784 10140 10836 10192
rect 13360 10208 13412 10260
rect 13452 10208 13504 10260
rect 22376 10251 22428 10260
rect 16304 10140 16356 10192
rect 11152 10115 11204 10124
rect 11152 10081 11161 10115
rect 11161 10081 11195 10115
rect 11195 10081 11204 10115
rect 11152 10072 11204 10081
rect 12256 10072 12308 10124
rect 5908 10004 5960 10056
rect 7104 10047 7156 10056
rect 5448 9979 5500 9988
rect 5448 9945 5482 9979
rect 5482 9945 5500 9979
rect 5448 9936 5500 9945
rect 7104 10013 7113 10047
rect 7113 10013 7147 10047
rect 7147 10013 7156 10047
rect 7104 10004 7156 10013
rect 8300 10004 8352 10056
rect 9220 10047 9272 10056
rect 9220 10013 9229 10047
rect 9229 10013 9263 10047
rect 9263 10013 9272 10047
rect 9220 10004 9272 10013
rect 9312 10047 9364 10056
rect 9312 10013 9321 10047
rect 9321 10013 9355 10047
rect 9355 10013 9364 10047
rect 12808 10047 12860 10056
rect 9312 10004 9364 10013
rect 12808 10013 12817 10047
rect 12817 10013 12851 10047
rect 12851 10013 12860 10047
rect 12808 10004 12860 10013
rect 13268 10004 13320 10056
rect 14188 10004 14240 10056
rect 15844 10072 15896 10124
rect 22376 10217 22385 10251
rect 22385 10217 22419 10251
rect 22419 10217 22428 10251
rect 22376 10208 22428 10217
rect 22560 10208 22612 10260
rect 17684 10183 17736 10192
rect 17684 10149 17693 10183
rect 17693 10149 17727 10183
rect 17727 10149 17736 10183
rect 17684 10140 17736 10149
rect 19248 10072 19300 10124
rect 14372 10004 14424 10056
rect 14740 10047 14792 10056
rect 14740 10013 14749 10047
rect 14749 10013 14783 10047
rect 14783 10013 14792 10047
rect 14740 10004 14792 10013
rect 15476 10004 15528 10056
rect 12072 9936 12124 9988
rect 13912 9936 13964 9988
rect 14004 9936 14056 9988
rect 14648 9936 14700 9988
rect 12348 9911 12400 9920
rect 12348 9877 12357 9911
rect 12357 9877 12391 9911
rect 12391 9877 12400 9911
rect 12348 9868 12400 9877
rect 14280 9911 14332 9920
rect 14280 9877 14289 9911
rect 14289 9877 14323 9911
rect 14323 9877 14332 9911
rect 14280 9868 14332 9877
rect 15384 9868 15436 9920
rect 15476 9868 15528 9920
rect 16764 10004 16816 10056
rect 18328 10047 18380 10056
rect 18328 10013 18337 10047
rect 18337 10013 18371 10047
rect 18371 10013 18380 10047
rect 18328 10004 18380 10013
rect 19156 10004 19208 10056
rect 19340 10047 19392 10056
rect 19340 10013 19349 10047
rect 19349 10013 19383 10047
rect 19383 10013 19392 10047
rect 19340 10004 19392 10013
rect 21916 10115 21968 10124
rect 21916 10081 21925 10115
rect 21925 10081 21959 10115
rect 21959 10081 21968 10115
rect 25688 10208 25740 10260
rect 21916 10072 21968 10081
rect 25504 10072 25556 10124
rect 22468 10004 22520 10056
rect 23480 10004 23532 10056
rect 23756 10004 23808 10056
rect 25780 10004 25832 10056
rect 27436 10047 27488 10056
rect 27436 10013 27445 10047
rect 27445 10013 27479 10047
rect 27479 10013 27488 10047
rect 27436 10004 27488 10013
rect 17592 9936 17644 9988
rect 16580 9868 16632 9920
rect 17960 9868 18012 9920
rect 21180 9911 21232 9920
rect 21180 9877 21189 9911
rect 21189 9877 21223 9911
rect 21223 9877 21232 9911
rect 21180 9868 21232 9877
rect 22008 9911 22060 9920
rect 22008 9877 22017 9911
rect 22017 9877 22051 9911
rect 22051 9877 22060 9911
rect 22008 9868 22060 9877
rect 23020 9936 23072 9988
rect 24492 9936 24544 9988
rect 24032 9911 24084 9920
rect 24032 9877 24041 9911
rect 24041 9877 24075 9911
rect 24075 9877 24084 9911
rect 24032 9868 24084 9877
rect 25136 9911 25188 9920
rect 25136 9877 25145 9911
rect 25145 9877 25179 9911
rect 25179 9877 25188 9911
rect 25136 9868 25188 9877
rect 10214 9766 10266 9818
rect 10278 9766 10330 9818
rect 10342 9766 10394 9818
rect 10406 9766 10458 9818
rect 10470 9766 10522 9818
rect 19478 9766 19530 9818
rect 19542 9766 19594 9818
rect 19606 9766 19658 9818
rect 19670 9766 19722 9818
rect 19734 9766 19786 9818
rect 7748 9596 7800 9648
rect 9128 9664 9180 9716
rect 14740 9707 14792 9716
rect 14740 9673 14749 9707
rect 14749 9673 14783 9707
rect 14783 9673 14792 9707
rect 14740 9664 14792 9673
rect 16764 9707 16816 9716
rect 16764 9673 16773 9707
rect 16773 9673 16807 9707
rect 16807 9673 16816 9707
rect 16764 9664 16816 9673
rect 20076 9664 20128 9716
rect 22008 9664 22060 9716
rect 22468 9664 22520 9716
rect 24032 9707 24084 9716
rect 8300 9639 8352 9648
rect 8300 9605 8309 9639
rect 8309 9605 8343 9639
rect 8343 9605 8352 9639
rect 8300 9596 8352 9605
rect 9312 9596 9364 9648
rect 11152 9596 11204 9648
rect 13084 9596 13136 9648
rect 17684 9596 17736 9648
rect 18144 9596 18196 9648
rect 21180 9596 21232 9648
rect 22560 9596 22612 9648
rect 24032 9673 24041 9707
rect 24041 9673 24075 9707
rect 24075 9673 24084 9707
rect 24032 9664 24084 9673
rect 24676 9707 24728 9716
rect 24676 9673 24685 9707
rect 24685 9673 24719 9707
rect 24719 9673 24728 9707
rect 24676 9664 24728 9673
rect 25136 9707 25188 9716
rect 25136 9673 25145 9707
rect 25145 9673 25179 9707
rect 25179 9673 25188 9707
rect 25136 9664 25188 9673
rect 26148 9664 26200 9716
rect 27436 9664 27488 9716
rect 24952 9596 25004 9648
rect 25688 9596 25740 9648
rect 26056 9639 26108 9648
rect 26056 9605 26065 9639
rect 26065 9605 26099 9639
rect 26099 9605 26108 9639
rect 26056 9596 26108 9605
rect 7380 9528 7432 9580
rect 8024 9571 8076 9580
rect 8024 9537 8033 9571
rect 8033 9537 8067 9571
rect 8067 9537 8076 9571
rect 8024 9528 8076 9537
rect 8668 9528 8720 9580
rect 9036 9571 9088 9580
rect 9036 9537 9045 9571
rect 9045 9537 9079 9571
rect 9079 9537 9088 9571
rect 9036 9528 9088 9537
rect 9128 9528 9180 9580
rect 9772 9571 9824 9580
rect 9772 9537 9806 9571
rect 9806 9537 9824 9571
rect 9772 9528 9824 9537
rect 12532 9571 12584 9580
rect 8852 9460 8904 9512
rect 8944 9460 8996 9512
rect 10508 9460 10560 9512
rect 12256 9460 12308 9512
rect 12532 9537 12541 9571
rect 12541 9537 12575 9571
rect 12575 9537 12584 9571
rect 12532 9528 12584 9537
rect 12716 9571 12768 9580
rect 12716 9537 12725 9571
rect 12725 9537 12759 9571
rect 12759 9537 12768 9571
rect 12716 9528 12768 9537
rect 12808 9571 12860 9580
rect 12808 9537 12817 9571
rect 12817 9537 12851 9571
rect 12851 9537 12860 9571
rect 12808 9528 12860 9537
rect 14464 9571 14516 9580
rect 14464 9537 14473 9571
rect 14473 9537 14507 9571
rect 14507 9537 14516 9571
rect 14464 9528 14516 9537
rect 15844 9528 15896 9580
rect 16304 9571 16356 9580
rect 14096 9503 14148 9512
rect 6920 9392 6972 9444
rect 14096 9469 14105 9503
rect 14105 9469 14139 9503
rect 14139 9469 14148 9503
rect 14096 9460 14148 9469
rect 16304 9537 16313 9571
rect 16313 9537 16347 9571
rect 16347 9537 16356 9571
rect 16304 9528 16356 9537
rect 17316 9571 17368 9580
rect 6000 9324 6052 9376
rect 7104 9324 7156 9376
rect 8024 9324 8076 9376
rect 8484 9367 8536 9376
rect 8484 9333 8493 9367
rect 8493 9333 8527 9367
rect 8527 9333 8536 9367
rect 8484 9324 8536 9333
rect 8668 9367 8720 9376
rect 8668 9333 8677 9367
rect 8677 9333 8711 9367
rect 8711 9333 8720 9367
rect 11152 9392 11204 9444
rect 12348 9392 12400 9444
rect 13728 9392 13780 9444
rect 16304 9392 16356 9444
rect 17316 9537 17325 9571
rect 17325 9537 17359 9571
rect 17359 9537 17368 9571
rect 17316 9528 17368 9537
rect 17408 9571 17460 9580
rect 17408 9537 17417 9571
rect 17417 9537 17451 9571
rect 17451 9537 17460 9571
rect 17408 9528 17460 9537
rect 17592 9571 17644 9580
rect 17592 9537 17601 9571
rect 17601 9537 17635 9571
rect 17635 9537 17644 9571
rect 18052 9571 18104 9580
rect 17592 9528 17644 9537
rect 18052 9537 18061 9571
rect 18061 9537 18095 9571
rect 18095 9537 18104 9571
rect 18052 9528 18104 9537
rect 10876 9367 10928 9376
rect 8668 9324 8720 9333
rect 10876 9333 10885 9367
rect 10885 9333 10919 9367
rect 10919 9333 10928 9367
rect 10876 9324 10928 9333
rect 11244 9324 11296 9376
rect 11428 9324 11480 9376
rect 12440 9324 12492 9376
rect 13636 9367 13688 9376
rect 13636 9333 13645 9367
rect 13645 9333 13679 9367
rect 13679 9333 13688 9367
rect 13636 9324 13688 9333
rect 17776 9324 17828 9376
rect 18236 9324 18288 9376
rect 21272 9571 21324 9580
rect 21272 9537 21281 9571
rect 21281 9537 21315 9571
rect 21315 9537 21324 9571
rect 21272 9528 21324 9537
rect 22192 9528 22244 9580
rect 23388 9528 23440 9580
rect 20536 9503 20588 9512
rect 20536 9469 20545 9503
rect 20545 9469 20579 9503
rect 20579 9469 20588 9503
rect 20536 9460 20588 9469
rect 24032 9392 24084 9444
rect 24860 9460 24912 9512
rect 24952 9392 25004 9444
rect 19708 9324 19760 9376
rect 23664 9367 23716 9376
rect 23664 9333 23673 9367
rect 23673 9333 23707 9367
rect 23707 9333 23716 9367
rect 23664 9324 23716 9333
rect 5582 9222 5634 9274
rect 5646 9222 5698 9274
rect 5710 9222 5762 9274
rect 5774 9222 5826 9274
rect 5838 9222 5890 9274
rect 14846 9222 14898 9274
rect 14910 9222 14962 9274
rect 14974 9222 15026 9274
rect 15038 9222 15090 9274
rect 15102 9222 15154 9274
rect 24110 9222 24162 9274
rect 24174 9222 24226 9274
rect 24238 9222 24290 9274
rect 24302 9222 24354 9274
rect 24366 9222 24418 9274
rect 7380 9163 7432 9172
rect 7380 9129 7389 9163
rect 7389 9129 7423 9163
rect 7423 9129 7432 9163
rect 7380 9120 7432 9129
rect 8484 9120 8536 9172
rect 9220 9120 9272 9172
rect 9772 9120 9824 9172
rect 8024 9052 8076 9104
rect 1860 8959 1912 8968
rect 1860 8925 1869 8959
rect 1869 8925 1903 8959
rect 1903 8925 1912 8959
rect 1860 8916 1912 8925
rect 4620 8916 4672 8968
rect 1676 8891 1728 8900
rect 1676 8857 1685 8891
rect 1685 8857 1719 8891
rect 1719 8857 1728 8891
rect 1676 8848 1728 8857
rect 6828 8848 6880 8900
rect 7932 8916 7984 8968
rect 8116 8959 8168 8968
rect 8116 8925 8125 8959
rect 8125 8925 8159 8959
rect 8159 8925 8168 8959
rect 10048 8984 10100 9036
rect 10508 8984 10560 9036
rect 13636 9120 13688 9172
rect 17316 9120 17368 9172
rect 10968 9052 11020 9104
rect 11520 9052 11572 9104
rect 15292 9095 15344 9104
rect 15292 9061 15301 9095
rect 15301 9061 15335 9095
rect 15335 9061 15344 9095
rect 15292 9052 15344 9061
rect 11428 8984 11480 9036
rect 11888 8984 11940 9036
rect 14004 8984 14056 9036
rect 8116 8916 8168 8925
rect 8392 8848 8444 8900
rect 8576 8848 8628 8900
rect 11428 8848 11480 8900
rect 11980 8916 12032 8968
rect 12440 8959 12492 8968
rect 12440 8925 12474 8959
rect 12474 8925 12492 8959
rect 12440 8916 12492 8925
rect 13636 8916 13688 8968
rect 15200 8984 15252 9036
rect 21272 9120 21324 9172
rect 20996 9052 21048 9104
rect 21732 9095 21784 9104
rect 21732 9061 21741 9095
rect 21741 9061 21775 9095
rect 21775 9061 21784 9095
rect 21732 9052 21784 9061
rect 22192 9120 22244 9172
rect 19708 9027 19760 9036
rect 19708 8993 19717 9027
rect 19717 8993 19751 9027
rect 19751 8993 19760 9027
rect 19708 8984 19760 8993
rect 7656 8823 7708 8832
rect 7656 8789 7665 8823
rect 7665 8789 7699 8823
rect 7699 8789 7708 8823
rect 7656 8780 7708 8789
rect 10140 8823 10192 8832
rect 10140 8789 10149 8823
rect 10149 8789 10183 8823
rect 10183 8789 10192 8823
rect 10140 8780 10192 8789
rect 13820 8848 13872 8900
rect 14464 8848 14516 8900
rect 15200 8848 15252 8900
rect 16672 8848 16724 8900
rect 17040 8848 17092 8900
rect 17592 8916 17644 8968
rect 17776 8959 17828 8968
rect 17776 8925 17810 8959
rect 17810 8925 17828 8959
rect 17776 8916 17828 8925
rect 18236 8916 18288 8968
rect 19892 8959 19944 8968
rect 19892 8925 19901 8959
rect 19901 8925 19935 8959
rect 19935 8925 19944 8959
rect 24860 8984 24912 9036
rect 19892 8916 19944 8925
rect 20720 8916 20772 8968
rect 21640 8959 21692 8968
rect 21640 8925 21649 8959
rect 21649 8925 21683 8959
rect 21683 8925 21692 8959
rect 21640 8916 21692 8925
rect 20444 8848 20496 8900
rect 22008 8916 22060 8968
rect 22836 8916 22888 8968
rect 12072 8780 12124 8832
rect 12256 8780 12308 8832
rect 12440 8780 12492 8832
rect 13084 8780 13136 8832
rect 17868 8780 17920 8832
rect 20536 8780 20588 8832
rect 21824 8780 21876 8832
rect 25136 8823 25188 8832
rect 25136 8789 25145 8823
rect 25145 8789 25179 8823
rect 25179 8789 25188 8823
rect 25136 8780 25188 8789
rect 25228 8823 25280 8832
rect 25228 8789 25237 8823
rect 25237 8789 25271 8823
rect 25271 8789 25280 8823
rect 28356 8959 28408 8968
rect 28356 8925 28365 8959
rect 28365 8925 28399 8959
rect 28399 8925 28408 8959
rect 28356 8916 28408 8925
rect 25228 8780 25280 8789
rect 25872 8823 25924 8832
rect 25872 8789 25881 8823
rect 25881 8789 25915 8823
rect 25915 8789 25924 8823
rect 25872 8780 25924 8789
rect 10214 8678 10266 8730
rect 10278 8678 10330 8730
rect 10342 8678 10394 8730
rect 10406 8678 10458 8730
rect 10470 8678 10522 8730
rect 19478 8678 19530 8730
rect 19542 8678 19594 8730
rect 19606 8678 19658 8730
rect 19670 8678 19722 8730
rect 19734 8678 19786 8730
rect 6828 8619 6880 8628
rect 6828 8585 6837 8619
rect 6837 8585 6871 8619
rect 6871 8585 6880 8619
rect 6828 8576 6880 8585
rect 8484 8576 8536 8628
rect 9496 8576 9548 8628
rect 10140 8576 10192 8628
rect 8576 8508 8628 8560
rect 1400 8440 1452 8492
rect 6368 8440 6420 8492
rect 7104 8483 7156 8492
rect 7104 8449 7113 8483
rect 7113 8449 7147 8483
rect 7147 8449 7156 8483
rect 7104 8440 7156 8449
rect 4620 8415 4672 8424
rect 4620 8381 4629 8415
rect 4629 8381 4663 8415
rect 4663 8381 4672 8415
rect 4620 8372 4672 8381
rect 7656 8372 7708 8424
rect 7932 8440 7984 8492
rect 8392 8483 8444 8492
rect 8392 8449 8401 8483
rect 8401 8449 8435 8483
rect 8435 8449 8444 8483
rect 8392 8440 8444 8449
rect 9680 8440 9732 8492
rect 10692 8508 10744 8560
rect 11428 8508 11480 8560
rect 12808 8576 12860 8628
rect 15844 8576 15896 8628
rect 17408 8576 17460 8628
rect 20076 8576 20128 8628
rect 20720 8576 20772 8628
rect 21640 8576 21692 8628
rect 25228 8576 25280 8628
rect 12440 8508 12492 8560
rect 12900 8508 12952 8560
rect 10416 8440 10468 8492
rect 10600 8440 10652 8492
rect 10876 8483 10928 8492
rect 10876 8449 10885 8483
rect 10885 8449 10919 8483
rect 10919 8449 10928 8483
rect 11520 8483 11572 8492
rect 10876 8440 10928 8449
rect 11520 8449 11529 8483
rect 11529 8449 11563 8483
rect 11563 8449 11572 8483
rect 11520 8440 11572 8449
rect 12072 8483 12124 8492
rect 12072 8449 12081 8483
rect 12081 8449 12115 8483
rect 12115 8449 12124 8483
rect 12072 8440 12124 8449
rect 13084 8483 13136 8492
rect 13084 8449 13093 8483
rect 13093 8449 13127 8483
rect 13127 8449 13136 8483
rect 13084 8440 13136 8449
rect 13268 8483 13320 8492
rect 13268 8449 13277 8483
rect 13277 8449 13311 8483
rect 13311 8449 13320 8483
rect 13268 8440 13320 8449
rect 14004 8440 14056 8492
rect 14280 8483 14332 8492
rect 14280 8449 14289 8483
rect 14289 8449 14323 8483
rect 14323 8449 14332 8483
rect 14280 8440 14332 8449
rect 14464 8483 14516 8492
rect 14464 8449 14473 8483
rect 14473 8449 14507 8483
rect 14507 8449 14516 8483
rect 14464 8440 14516 8449
rect 16212 8508 16264 8560
rect 17040 8508 17092 8560
rect 15200 8483 15252 8492
rect 15200 8449 15234 8483
rect 15234 8449 15252 8483
rect 15200 8440 15252 8449
rect 17868 8508 17920 8560
rect 19156 8551 19208 8560
rect 19156 8517 19165 8551
rect 19165 8517 19199 8551
rect 19199 8517 19208 8551
rect 19156 8508 19208 8517
rect 19432 8508 19484 8560
rect 19892 8508 19944 8560
rect 22652 8551 22704 8560
rect 22652 8517 22661 8551
rect 22661 8517 22695 8551
rect 22695 8517 22704 8551
rect 22652 8508 22704 8517
rect 22836 8551 22888 8560
rect 22836 8517 22845 8551
rect 22845 8517 22879 8551
rect 22879 8517 22888 8551
rect 22836 8508 22888 8517
rect 19984 8483 20036 8492
rect 19984 8449 20018 8483
rect 20018 8449 20036 8483
rect 10692 8372 10744 8424
rect 11796 8415 11848 8424
rect 6092 8236 6144 8288
rect 6920 8236 6972 8288
rect 7656 8279 7708 8288
rect 7656 8245 7665 8279
rect 7665 8245 7699 8279
rect 7699 8245 7708 8279
rect 7656 8236 7708 8245
rect 10508 8304 10560 8356
rect 11796 8381 11805 8415
rect 11805 8381 11839 8415
rect 11839 8381 11848 8415
rect 11796 8372 11848 8381
rect 11888 8372 11940 8424
rect 12256 8372 12308 8424
rect 14096 8372 14148 8424
rect 14740 8372 14792 8424
rect 19984 8440 20036 8449
rect 23756 8483 23808 8492
rect 23756 8449 23790 8483
rect 23790 8449 23808 8483
rect 25872 8508 25924 8560
rect 23756 8440 23808 8449
rect 12348 8347 12400 8356
rect 10692 8236 10744 8288
rect 12348 8313 12357 8347
rect 12357 8313 12391 8347
rect 12391 8313 12400 8347
rect 12348 8304 12400 8313
rect 16948 8304 17000 8356
rect 17592 8372 17644 8424
rect 23480 8415 23532 8424
rect 18696 8347 18748 8356
rect 18696 8313 18705 8347
rect 18705 8313 18739 8347
rect 18739 8313 18748 8347
rect 18696 8304 18748 8313
rect 19340 8304 19392 8356
rect 11244 8236 11296 8288
rect 11612 8279 11664 8288
rect 11612 8245 11621 8279
rect 11621 8245 11655 8279
rect 11655 8245 11664 8279
rect 11612 8236 11664 8245
rect 13176 8279 13228 8288
rect 13176 8245 13185 8279
rect 13185 8245 13219 8279
rect 13219 8245 13228 8279
rect 13176 8236 13228 8245
rect 14188 8236 14240 8288
rect 14464 8236 14516 8288
rect 15568 8236 15620 8288
rect 23480 8381 23489 8415
rect 23489 8381 23523 8415
rect 23523 8381 23532 8415
rect 23480 8372 23532 8381
rect 21088 8347 21140 8356
rect 21088 8313 21097 8347
rect 21097 8313 21131 8347
rect 21131 8313 21140 8347
rect 21088 8304 21140 8313
rect 19892 8236 19944 8288
rect 26148 8236 26200 8288
rect 5582 8134 5634 8186
rect 5646 8134 5698 8186
rect 5710 8134 5762 8186
rect 5774 8134 5826 8186
rect 5838 8134 5890 8186
rect 14846 8134 14898 8186
rect 14910 8134 14962 8186
rect 14974 8134 15026 8186
rect 15038 8134 15090 8186
rect 15102 8134 15154 8186
rect 24110 8134 24162 8186
rect 24174 8134 24226 8186
rect 24238 8134 24290 8186
rect 24302 8134 24354 8186
rect 24366 8134 24418 8186
rect 1400 8075 1452 8084
rect 1400 8041 1409 8075
rect 1409 8041 1443 8075
rect 1443 8041 1452 8075
rect 1400 8032 1452 8041
rect 6368 8075 6420 8084
rect 6368 8041 6377 8075
rect 6377 8041 6411 8075
rect 6411 8041 6420 8075
rect 6368 8032 6420 8041
rect 10416 8032 10468 8084
rect 10876 8032 10928 8084
rect 11520 8075 11572 8084
rect 11520 8041 11529 8075
rect 11529 8041 11563 8075
rect 11563 8041 11572 8075
rect 11520 8032 11572 8041
rect 12072 8032 12124 8084
rect 12716 8032 12768 8084
rect 12900 8032 12952 8084
rect 14188 8032 14240 8084
rect 15200 8032 15252 8084
rect 15292 8032 15344 8084
rect 16212 8075 16264 8084
rect 16212 8041 16221 8075
rect 16221 8041 16255 8075
rect 16255 8041 16264 8075
rect 16212 8032 16264 8041
rect 16488 8075 16540 8084
rect 16488 8041 16497 8075
rect 16497 8041 16531 8075
rect 16531 8041 16540 8075
rect 16488 8032 16540 8041
rect 16948 8075 17000 8084
rect 16948 8041 16957 8075
rect 16957 8041 16991 8075
rect 16991 8041 17000 8075
rect 16948 8032 17000 8041
rect 18052 8032 18104 8084
rect 18328 8032 18380 8084
rect 18512 8032 18564 8084
rect 19984 8032 20036 8084
rect 7012 7964 7064 8016
rect 6092 7939 6144 7948
rect 6092 7905 6101 7939
rect 6101 7905 6135 7939
rect 6135 7905 6144 7939
rect 6092 7896 6144 7905
rect 5908 7871 5960 7880
rect 5908 7837 5917 7871
rect 5917 7837 5951 7871
rect 5951 7837 5960 7871
rect 10508 7939 10560 7948
rect 10508 7905 10517 7939
rect 10517 7905 10551 7939
rect 10551 7905 10560 7939
rect 10508 7896 10560 7905
rect 5908 7828 5960 7837
rect 6920 7828 6972 7880
rect 7012 7871 7064 7880
rect 7012 7837 7021 7871
rect 7021 7837 7055 7871
rect 7055 7837 7064 7871
rect 7564 7871 7616 7880
rect 7012 7828 7064 7837
rect 7564 7837 7573 7871
rect 7573 7837 7607 7871
rect 7607 7837 7616 7871
rect 7564 7828 7616 7837
rect 7840 7828 7892 7880
rect 8024 7871 8076 7880
rect 8024 7837 8033 7871
rect 8033 7837 8067 7871
rect 8067 7837 8076 7871
rect 8024 7828 8076 7837
rect 10048 7871 10100 7880
rect 6460 7760 6512 7812
rect 6644 7803 6696 7812
rect 6644 7769 6653 7803
rect 6653 7769 6687 7803
rect 6687 7769 6696 7803
rect 6644 7760 6696 7769
rect 6736 7803 6788 7812
rect 6736 7769 6745 7803
rect 6745 7769 6779 7803
rect 6779 7769 6788 7803
rect 10048 7837 10057 7871
rect 10057 7837 10091 7871
rect 10091 7837 10100 7871
rect 10048 7828 10100 7837
rect 10600 7828 10652 7880
rect 12440 7896 12492 7948
rect 6736 7760 6788 7769
rect 7840 7692 7892 7744
rect 11060 7760 11112 7812
rect 10692 7692 10744 7744
rect 11796 7871 11848 7880
rect 11796 7837 11805 7871
rect 11805 7837 11839 7871
rect 11839 7837 11848 7871
rect 11796 7828 11848 7837
rect 12256 7871 12308 7880
rect 12256 7837 12265 7871
rect 12265 7837 12299 7871
rect 12299 7837 12308 7871
rect 12256 7828 12308 7837
rect 11612 7760 11664 7812
rect 13084 7896 13136 7948
rect 13360 7896 13412 7948
rect 15568 7939 15620 7948
rect 13268 7828 13320 7880
rect 15568 7905 15577 7939
rect 15577 7905 15611 7939
rect 15611 7905 15620 7939
rect 15568 7896 15620 7905
rect 18604 7964 18656 8016
rect 19616 7964 19668 8016
rect 20628 8032 20680 8084
rect 22284 8032 22336 8084
rect 23756 8075 23808 8084
rect 23756 8041 23765 8075
rect 23765 8041 23799 8075
rect 23799 8041 23808 8075
rect 23756 8032 23808 8041
rect 25136 8032 25188 8084
rect 20536 7964 20588 8016
rect 21732 7964 21784 8016
rect 19156 7896 19208 7948
rect 19340 7939 19392 7948
rect 19340 7905 19349 7939
rect 19349 7905 19383 7939
rect 19383 7905 19392 7939
rect 19340 7896 19392 7905
rect 25872 7939 25924 7948
rect 13636 7760 13688 7812
rect 14280 7803 14332 7812
rect 14280 7769 14307 7803
rect 14307 7769 14332 7803
rect 14280 7760 14332 7769
rect 17040 7871 17092 7880
rect 17040 7837 17049 7871
rect 17049 7837 17083 7871
rect 17083 7837 17092 7871
rect 17040 7828 17092 7837
rect 17868 7828 17920 7880
rect 18328 7828 18380 7880
rect 19616 7828 19668 7880
rect 19984 7828 20036 7880
rect 20444 7871 20496 7880
rect 20444 7837 20453 7871
rect 20453 7837 20487 7871
rect 20487 7837 20496 7871
rect 20444 7828 20496 7837
rect 20536 7871 20588 7880
rect 20536 7837 20545 7871
rect 20545 7837 20579 7871
rect 20579 7837 20588 7871
rect 20536 7828 20588 7837
rect 20996 7828 21048 7880
rect 16488 7692 16540 7744
rect 20628 7760 20680 7812
rect 25872 7905 25881 7939
rect 25881 7905 25915 7939
rect 25915 7905 25924 7939
rect 25872 7896 25924 7905
rect 17316 7735 17368 7744
rect 17316 7701 17325 7735
rect 17325 7701 17359 7735
rect 17359 7701 17368 7735
rect 17316 7692 17368 7701
rect 18512 7692 18564 7744
rect 20260 7692 20312 7744
rect 20904 7735 20956 7744
rect 20904 7701 20913 7735
rect 20913 7701 20947 7735
rect 20947 7701 20956 7735
rect 20904 7692 20956 7701
rect 21180 7692 21232 7744
rect 23480 7828 23532 7880
rect 23664 7828 23716 7880
rect 23940 7828 23992 7880
rect 25412 7828 25464 7880
rect 26148 7828 26200 7880
rect 28356 7871 28408 7880
rect 28356 7837 28365 7871
rect 28365 7837 28399 7871
rect 28399 7837 28408 7871
rect 28356 7828 28408 7837
rect 21364 7692 21416 7744
rect 22652 7692 22704 7744
rect 25780 7692 25832 7744
rect 10214 7590 10266 7642
rect 10278 7590 10330 7642
rect 10342 7590 10394 7642
rect 10406 7590 10458 7642
rect 10470 7590 10522 7642
rect 19478 7590 19530 7642
rect 19542 7590 19594 7642
rect 19606 7590 19658 7642
rect 19670 7590 19722 7642
rect 19734 7590 19786 7642
rect 8116 7488 8168 7540
rect 10968 7488 11020 7540
rect 11888 7488 11940 7540
rect 14464 7488 14516 7540
rect 17408 7531 17460 7540
rect 7840 7463 7892 7472
rect 7840 7429 7849 7463
rect 7849 7429 7883 7463
rect 7883 7429 7892 7463
rect 7840 7420 7892 7429
rect 11060 7420 11112 7472
rect 4620 7395 4672 7404
rect 4620 7361 4629 7395
rect 4629 7361 4663 7395
rect 4663 7361 4672 7395
rect 4620 7352 4672 7361
rect 7012 7352 7064 7404
rect 7656 7395 7708 7404
rect 7656 7361 7665 7395
rect 7665 7361 7699 7395
rect 7699 7361 7708 7395
rect 7656 7352 7708 7361
rect 6460 7284 6512 7336
rect 7564 7284 7616 7336
rect 8484 7352 8536 7404
rect 9128 7259 9180 7268
rect 9128 7225 9137 7259
rect 9137 7225 9171 7259
rect 9171 7225 9180 7259
rect 9128 7216 9180 7225
rect 9864 7352 9916 7404
rect 10508 7352 10560 7404
rect 11152 7352 11204 7404
rect 11520 7352 11572 7404
rect 10784 7284 10836 7336
rect 13268 7420 13320 7472
rect 17408 7497 17417 7531
rect 17417 7497 17451 7531
rect 17451 7497 17460 7531
rect 17408 7488 17460 7497
rect 17500 7488 17552 7540
rect 20904 7488 20956 7540
rect 12440 7352 12492 7404
rect 12624 7352 12676 7404
rect 14372 7352 14424 7404
rect 15476 7420 15528 7472
rect 16488 7420 16540 7472
rect 15844 7395 15896 7404
rect 12164 7284 12216 7336
rect 9772 7216 9824 7268
rect 13176 7284 13228 7336
rect 14648 7284 14700 7336
rect 15844 7361 15853 7395
rect 15853 7361 15887 7395
rect 15887 7361 15896 7395
rect 15844 7352 15896 7361
rect 15936 7395 15988 7404
rect 15936 7361 15945 7395
rect 15945 7361 15979 7395
rect 15979 7361 15988 7395
rect 15936 7352 15988 7361
rect 17040 7352 17092 7404
rect 19984 7420 20036 7472
rect 20536 7420 20588 7472
rect 20996 7463 21048 7472
rect 20996 7429 21005 7463
rect 21005 7429 21039 7463
rect 21039 7429 21048 7463
rect 20996 7420 21048 7429
rect 21180 7420 21232 7472
rect 21824 7463 21876 7472
rect 21824 7429 21833 7463
rect 21833 7429 21867 7463
rect 21867 7429 21876 7463
rect 21824 7420 21876 7429
rect 24032 7488 24084 7540
rect 25228 7488 25280 7540
rect 22652 7463 22704 7472
rect 22652 7429 22661 7463
rect 22661 7429 22695 7463
rect 22695 7429 22704 7463
rect 22652 7420 22704 7429
rect 24492 7463 24544 7472
rect 17500 7395 17552 7404
rect 17500 7361 17509 7395
rect 17509 7361 17543 7395
rect 17543 7361 17552 7395
rect 17500 7352 17552 7361
rect 17592 7352 17644 7404
rect 19340 7352 19392 7404
rect 19708 7352 19760 7404
rect 20812 7395 20864 7404
rect 20812 7361 20821 7395
rect 20821 7361 20855 7395
rect 20855 7361 20864 7395
rect 20812 7352 20864 7361
rect 12900 7216 12952 7268
rect 19984 7284 20036 7336
rect 21640 7284 21692 7336
rect 24492 7429 24501 7463
rect 24501 7429 24535 7463
rect 24535 7429 24544 7463
rect 24492 7420 24544 7429
rect 24952 7420 25004 7472
rect 24860 7352 24912 7404
rect 21364 7216 21416 7268
rect 22284 7327 22336 7336
rect 22284 7293 22293 7327
rect 22293 7293 22327 7327
rect 22327 7293 22336 7327
rect 22284 7284 22336 7293
rect 22836 7284 22888 7336
rect 25872 7284 25924 7336
rect 23572 7259 23624 7268
rect 23572 7225 23581 7259
rect 23581 7225 23615 7259
rect 23615 7225 23624 7259
rect 23572 7216 23624 7225
rect 9864 7191 9916 7200
rect 9864 7157 9873 7191
rect 9873 7157 9907 7191
rect 9907 7157 9916 7191
rect 9864 7148 9916 7157
rect 9956 7148 10008 7200
rect 11612 7148 11664 7200
rect 14372 7148 14424 7200
rect 16028 7148 16080 7200
rect 18420 7148 18472 7200
rect 19064 7148 19116 7200
rect 21732 7148 21784 7200
rect 22836 7191 22888 7200
rect 22836 7157 22845 7191
rect 22845 7157 22879 7191
rect 22879 7157 22888 7191
rect 22836 7148 22888 7157
rect 23112 7148 23164 7200
rect 25320 7148 25372 7200
rect 5582 7046 5634 7098
rect 5646 7046 5698 7098
rect 5710 7046 5762 7098
rect 5774 7046 5826 7098
rect 5838 7046 5890 7098
rect 14846 7046 14898 7098
rect 14910 7046 14962 7098
rect 14974 7046 15026 7098
rect 15038 7046 15090 7098
rect 15102 7046 15154 7098
rect 24110 7046 24162 7098
rect 24174 7046 24226 7098
rect 24238 7046 24290 7098
rect 24302 7046 24354 7098
rect 24366 7046 24418 7098
rect 5908 6944 5960 6996
rect 7104 6944 7156 6996
rect 8024 6944 8076 6996
rect 8392 6944 8444 6996
rect 8576 6944 8628 6996
rect 4620 6876 4672 6928
rect 7932 6876 7984 6928
rect 6920 6783 6972 6792
rect 6920 6749 6929 6783
rect 6929 6749 6963 6783
rect 6963 6749 6972 6783
rect 6920 6740 6972 6749
rect 7012 6783 7064 6792
rect 7012 6749 7021 6783
rect 7021 6749 7055 6783
rect 7055 6749 7064 6783
rect 7932 6783 7984 6792
rect 7012 6740 7064 6749
rect 7932 6749 7941 6783
rect 7941 6749 7975 6783
rect 7975 6749 7984 6783
rect 7932 6740 7984 6749
rect 6368 6715 6420 6724
rect 6368 6681 6386 6715
rect 6386 6681 6420 6715
rect 6368 6672 6420 6681
rect 5908 6604 5960 6656
rect 7748 6647 7800 6656
rect 7748 6613 7757 6647
rect 7757 6613 7791 6647
rect 7791 6613 7800 6647
rect 7748 6604 7800 6613
rect 8392 6740 8444 6792
rect 9128 6944 9180 6996
rect 9220 6944 9272 6996
rect 10508 6944 10560 6996
rect 12532 6944 12584 6996
rect 15476 6987 15528 6996
rect 15476 6953 15485 6987
rect 15485 6953 15519 6987
rect 15519 6953 15528 6987
rect 15476 6944 15528 6953
rect 17408 6944 17460 6996
rect 18420 6987 18472 6996
rect 18420 6953 18429 6987
rect 18429 6953 18463 6987
rect 18463 6953 18472 6987
rect 18420 6944 18472 6953
rect 20536 6987 20588 6996
rect 20536 6953 20545 6987
rect 20545 6953 20579 6987
rect 20579 6953 20588 6987
rect 20536 6944 20588 6953
rect 23940 6944 23992 6996
rect 12164 6919 12216 6928
rect 12164 6885 12173 6919
rect 12173 6885 12207 6919
rect 12207 6885 12216 6919
rect 12164 6876 12216 6885
rect 10784 6783 10836 6792
rect 8300 6604 8352 6656
rect 9680 6672 9732 6724
rect 10784 6749 10793 6783
rect 10793 6749 10827 6783
rect 10827 6749 10836 6783
rect 10784 6740 10836 6749
rect 11888 6808 11940 6860
rect 17500 6876 17552 6928
rect 11152 6783 11204 6792
rect 11152 6749 11161 6783
rect 11161 6749 11195 6783
rect 11195 6749 11204 6783
rect 11152 6740 11204 6749
rect 11336 6740 11388 6792
rect 11704 6740 11756 6792
rect 10048 6604 10100 6656
rect 10600 6647 10652 6656
rect 10600 6613 10609 6647
rect 10609 6613 10643 6647
rect 10643 6613 10652 6647
rect 10600 6604 10652 6613
rect 11428 6672 11480 6724
rect 17316 6808 17368 6860
rect 11336 6604 11388 6656
rect 11796 6604 11848 6656
rect 12716 6740 12768 6792
rect 12900 6783 12952 6792
rect 12900 6749 12909 6783
rect 12909 6749 12943 6783
rect 12943 6749 12952 6783
rect 12900 6740 12952 6749
rect 13636 6783 13688 6792
rect 13636 6749 13645 6783
rect 13645 6749 13679 6783
rect 13679 6749 13688 6783
rect 13636 6740 13688 6749
rect 13912 6740 13964 6792
rect 14740 6740 14792 6792
rect 16028 6783 16080 6792
rect 16028 6749 16062 6783
rect 16062 6749 16080 6783
rect 16028 6740 16080 6749
rect 24952 6919 25004 6928
rect 14188 6672 14240 6724
rect 17776 6740 17828 6792
rect 24952 6885 24961 6919
rect 24961 6885 24995 6919
rect 24995 6885 25004 6919
rect 24952 6876 25004 6885
rect 18696 6783 18748 6792
rect 18696 6749 18705 6783
rect 18705 6749 18739 6783
rect 18739 6749 18748 6783
rect 18696 6740 18748 6749
rect 19248 6783 19300 6792
rect 19248 6749 19257 6783
rect 19257 6749 19291 6783
rect 19291 6749 19300 6783
rect 19248 6740 19300 6749
rect 19524 6740 19576 6792
rect 20444 6808 20496 6860
rect 22100 6808 22152 6860
rect 20812 6740 20864 6792
rect 21088 6783 21140 6792
rect 21088 6749 21097 6783
rect 21097 6749 21131 6783
rect 21131 6749 21140 6783
rect 21088 6740 21140 6749
rect 21272 6783 21324 6792
rect 21272 6749 21281 6783
rect 21281 6749 21315 6783
rect 21315 6749 21324 6783
rect 21272 6740 21324 6749
rect 19708 6715 19760 6724
rect 19708 6681 19717 6715
rect 19717 6681 19751 6715
rect 19751 6681 19760 6715
rect 19708 6672 19760 6681
rect 21640 6715 21692 6724
rect 12440 6604 12492 6656
rect 12808 6647 12860 6656
rect 12808 6613 12817 6647
rect 12817 6613 12851 6647
rect 12851 6613 12860 6647
rect 12808 6604 12860 6613
rect 14004 6604 14056 6656
rect 17132 6647 17184 6656
rect 17132 6613 17141 6647
rect 17141 6613 17175 6647
rect 17175 6613 17184 6647
rect 17132 6604 17184 6613
rect 17500 6604 17552 6656
rect 19984 6604 20036 6656
rect 21640 6681 21649 6715
rect 21649 6681 21683 6715
rect 21683 6681 21692 6715
rect 21640 6672 21692 6681
rect 22008 6672 22060 6724
rect 22928 6715 22980 6724
rect 22928 6681 22962 6715
rect 22962 6681 22980 6715
rect 22928 6672 22980 6681
rect 23572 6672 23624 6724
rect 24676 6672 24728 6724
rect 25688 6672 25740 6724
rect 23388 6604 23440 6656
rect 25136 6604 25188 6656
rect 10214 6502 10266 6554
rect 10278 6502 10330 6554
rect 10342 6502 10394 6554
rect 10406 6502 10458 6554
rect 10470 6502 10522 6554
rect 19478 6502 19530 6554
rect 19542 6502 19594 6554
rect 19606 6502 19658 6554
rect 19670 6502 19722 6554
rect 19734 6502 19786 6554
rect 6368 6400 6420 6452
rect 6644 6400 6696 6452
rect 8116 6400 8168 6452
rect 8392 6443 8444 6452
rect 8392 6409 8401 6443
rect 8401 6409 8435 6443
rect 8435 6409 8444 6443
rect 8392 6400 8444 6409
rect 8484 6400 8536 6452
rect 9864 6443 9916 6452
rect 9864 6409 9873 6443
rect 9873 6409 9907 6443
rect 9907 6409 9916 6443
rect 9864 6400 9916 6409
rect 9956 6400 10008 6452
rect 12716 6400 12768 6452
rect 14188 6443 14240 6452
rect 14188 6409 14203 6443
rect 14203 6409 14237 6443
rect 14237 6409 14240 6443
rect 14188 6400 14240 6409
rect 15936 6400 15988 6452
rect 7748 6332 7800 6384
rect 6828 6307 6880 6316
rect 6828 6273 6837 6307
rect 6837 6273 6871 6307
rect 6871 6273 6880 6307
rect 7104 6307 7156 6316
rect 6828 6264 6880 6273
rect 7104 6273 7113 6307
rect 7113 6273 7147 6307
rect 7147 6273 7156 6307
rect 7104 6264 7156 6273
rect 7564 6307 7616 6316
rect 7564 6273 7573 6307
rect 7573 6273 7607 6307
rect 7607 6273 7616 6307
rect 7564 6264 7616 6273
rect 9772 6332 9824 6384
rect 8300 6196 8352 6248
rect 10600 6264 10652 6316
rect 11060 6332 11112 6384
rect 9864 6196 9916 6248
rect 10140 6196 10192 6248
rect 11888 6196 11940 6248
rect 13912 6332 13964 6384
rect 14648 6332 14700 6384
rect 12256 6264 12308 6316
rect 14004 6264 14056 6316
rect 14372 6307 14424 6316
rect 14372 6273 14381 6307
rect 14381 6273 14415 6307
rect 14415 6273 14424 6307
rect 14372 6264 14424 6273
rect 15476 6264 15528 6316
rect 17500 6264 17552 6316
rect 17132 6196 17184 6248
rect 17960 6400 18012 6452
rect 18696 6400 18748 6452
rect 18052 6332 18104 6384
rect 18604 6332 18656 6384
rect 21272 6400 21324 6452
rect 18972 6264 19024 6316
rect 20260 6375 20312 6384
rect 20260 6341 20269 6375
rect 20269 6341 20303 6375
rect 20303 6341 20312 6375
rect 20260 6332 20312 6341
rect 8484 6128 8536 6180
rect 9680 6171 9732 6180
rect 9680 6137 9689 6171
rect 9689 6137 9723 6171
rect 9723 6137 9732 6171
rect 9680 6128 9732 6137
rect 11980 6128 12032 6180
rect 7564 6060 7616 6112
rect 12072 6060 12124 6112
rect 12348 6060 12400 6112
rect 17776 6196 17828 6248
rect 19984 6264 20036 6316
rect 21088 6264 21140 6316
rect 21364 6196 21416 6248
rect 22928 6375 22980 6384
rect 22928 6341 22937 6375
rect 22937 6341 22971 6375
rect 22971 6341 22980 6375
rect 22928 6332 22980 6341
rect 22008 6264 22060 6316
rect 23112 6307 23164 6316
rect 23112 6273 23121 6307
rect 23121 6273 23155 6307
rect 23155 6273 23164 6307
rect 23112 6264 23164 6273
rect 17408 6128 17460 6180
rect 19432 6128 19484 6180
rect 20076 6128 20128 6180
rect 20996 6128 21048 6180
rect 23020 6239 23072 6248
rect 23020 6205 23029 6239
rect 23029 6205 23063 6239
rect 23063 6205 23072 6239
rect 23020 6196 23072 6205
rect 17868 6060 17920 6112
rect 19064 6103 19116 6112
rect 19064 6069 19073 6103
rect 19073 6069 19107 6103
rect 19107 6069 19116 6103
rect 19064 6060 19116 6069
rect 20260 6060 20312 6112
rect 21824 6060 21876 6112
rect 22192 6060 22244 6112
rect 23940 6400 23992 6452
rect 25688 6443 25740 6452
rect 25688 6409 25697 6443
rect 25697 6409 25731 6443
rect 25731 6409 25740 6443
rect 25688 6400 25740 6409
rect 25320 6375 25372 6384
rect 25320 6341 25329 6375
rect 25329 6341 25363 6375
rect 25363 6341 25372 6375
rect 25320 6332 25372 6341
rect 25412 6375 25464 6384
rect 25412 6341 25421 6375
rect 25421 6341 25455 6375
rect 25455 6341 25464 6375
rect 25412 6332 25464 6341
rect 23388 6307 23440 6316
rect 23388 6273 23397 6307
rect 23397 6273 23431 6307
rect 23431 6273 23440 6307
rect 23848 6307 23900 6316
rect 23388 6264 23440 6273
rect 23848 6273 23857 6307
rect 23857 6273 23891 6307
rect 23891 6273 23900 6307
rect 23848 6264 23900 6273
rect 24676 6307 24728 6316
rect 24676 6273 24685 6307
rect 24685 6273 24719 6307
rect 24719 6273 24728 6307
rect 24676 6264 24728 6273
rect 25136 6307 25188 6316
rect 25136 6273 25145 6307
rect 25145 6273 25179 6307
rect 25179 6273 25188 6307
rect 25136 6264 25188 6273
rect 24860 6171 24912 6180
rect 24860 6137 24869 6171
rect 24869 6137 24903 6171
rect 24903 6137 24912 6171
rect 24860 6128 24912 6137
rect 24032 6103 24084 6112
rect 24032 6069 24041 6103
rect 24041 6069 24075 6103
rect 24075 6069 24084 6103
rect 24032 6060 24084 6069
rect 5582 5958 5634 6010
rect 5646 5958 5698 6010
rect 5710 5958 5762 6010
rect 5774 5958 5826 6010
rect 5838 5958 5890 6010
rect 14846 5958 14898 6010
rect 14910 5958 14962 6010
rect 14974 5958 15026 6010
rect 15038 5958 15090 6010
rect 15102 5958 15154 6010
rect 24110 5958 24162 6010
rect 24174 5958 24226 6010
rect 24238 5958 24290 6010
rect 24302 5958 24354 6010
rect 24366 5958 24418 6010
rect 8484 5899 8536 5908
rect 8484 5865 8493 5899
rect 8493 5865 8527 5899
rect 8527 5865 8536 5899
rect 8484 5856 8536 5865
rect 10692 5856 10744 5908
rect 12256 5856 12308 5908
rect 12900 5856 12952 5908
rect 13360 5856 13412 5908
rect 8116 5763 8168 5772
rect 8116 5729 8125 5763
rect 8125 5729 8159 5763
rect 8159 5729 8168 5763
rect 8116 5720 8168 5729
rect 8576 5720 8628 5772
rect 1492 5559 1544 5568
rect 1492 5525 1501 5559
rect 1501 5525 1535 5559
rect 1535 5525 1544 5559
rect 1492 5516 1544 5525
rect 8484 5652 8536 5704
rect 9680 5788 9732 5840
rect 9312 5763 9364 5772
rect 9312 5729 9321 5763
rect 9321 5729 9355 5763
rect 9355 5729 9364 5763
rect 9312 5720 9364 5729
rect 12348 5788 12400 5840
rect 12532 5788 12584 5840
rect 12716 5788 12768 5840
rect 19064 5856 19116 5908
rect 19432 5899 19484 5908
rect 19432 5865 19441 5899
rect 19441 5865 19475 5899
rect 19475 5865 19484 5899
rect 19432 5856 19484 5865
rect 21272 5856 21324 5908
rect 22192 5899 22244 5908
rect 22192 5865 22201 5899
rect 22201 5865 22235 5899
rect 22235 5865 22244 5899
rect 22192 5856 22244 5865
rect 15384 5788 15436 5840
rect 16948 5788 17000 5840
rect 10784 5720 10836 5772
rect 9588 5559 9640 5568
rect 9588 5525 9597 5559
rect 9597 5525 9631 5559
rect 9631 5525 9640 5559
rect 9588 5516 9640 5525
rect 10048 5695 10100 5704
rect 10048 5661 10057 5695
rect 10057 5661 10091 5695
rect 10091 5661 10100 5695
rect 10048 5652 10100 5661
rect 10140 5695 10192 5704
rect 10140 5661 10149 5695
rect 10149 5661 10183 5695
rect 10183 5661 10192 5695
rect 10140 5652 10192 5661
rect 10600 5652 10652 5704
rect 13176 5720 13228 5772
rect 11520 5695 11572 5704
rect 11060 5584 11112 5636
rect 11520 5661 11529 5695
rect 11529 5661 11563 5695
rect 11563 5661 11572 5695
rect 11520 5652 11572 5661
rect 11704 5695 11756 5704
rect 11704 5661 11713 5695
rect 11713 5661 11747 5695
rect 11747 5661 11756 5695
rect 11704 5652 11756 5661
rect 11796 5695 11848 5704
rect 11796 5661 11805 5695
rect 11805 5661 11839 5695
rect 11839 5661 11848 5695
rect 11796 5652 11848 5661
rect 12072 5652 12124 5704
rect 12440 5652 12492 5704
rect 13912 5652 13964 5704
rect 16580 5695 16632 5704
rect 16580 5661 16589 5695
rect 16589 5661 16623 5695
rect 16623 5661 16632 5695
rect 16580 5652 16632 5661
rect 18788 5788 18840 5840
rect 17776 5720 17828 5772
rect 21824 5788 21876 5840
rect 12164 5584 12216 5636
rect 9956 5516 10008 5568
rect 10692 5559 10744 5568
rect 10692 5525 10701 5559
rect 10701 5525 10735 5559
rect 10735 5525 10744 5559
rect 10692 5516 10744 5525
rect 11336 5516 11388 5568
rect 11796 5516 11848 5568
rect 13084 5584 13136 5636
rect 13360 5584 13412 5636
rect 14556 5627 14608 5636
rect 14556 5593 14565 5627
rect 14565 5593 14599 5627
rect 14599 5593 14608 5627
rect 14556 5584 14608 5593
rect 17868 5652 17920 5704
rect 17960 5652 18012 5704
rect 18328 5695 18380 5704
rect 18328 5661 18337 5695
rect 18337 5661 18371 5695
rect 18371 5661 18380 5695
rect 18328 5652 18380 5661
rect 19892 5720 19944 5772
rect 20996 5720 21048 5772
rect 23848 5856 23900 5908
rect 23756 5788 23808 5840
rect 24676 5720 24728 5772
rect 20260 5695 20312 5704
rect 20260 5661 20294 5695
rect 20294 5661 20312 5695
rect 20260 5652 20312 5661
rect 21364 5652 21416 5704
rect 22100 5652 22152 5704
rect 18144 5584 18196 5636
rect 14280 5516 14332 5568
rect 17408 5516 17460 5568
rect 17868 5516 17920 5568
rect 19340 5584 19392 5636
rect 22652 5695 22704 5704
rect 22652 5661 22661 5695
rect 22661 5661 22695 5695
rect 22695 5661 22704 5695
rect 22652 5652 22704 5661
rect 23756 5695 23808 5704
rect 23756 5661 23765 5695
rect 23765 5661 23799 5695
rect 23799 5661 23808 5695
rect 23756 5652 23808 5661
rect 25136 5652 25188 5704
rect 28356 5695 28408 5704
rect 28356 5661 28365 5695
rect 28365 5661 28399 5695
rect 28399 5661 28408 5695
rect 28356 5652 28408 5661
rect 18972 5516 19024 5568
rect 20352 5516 20404 5568
rect 22560 5516 22612 5568
rect 23020 5516 23072 5568
rect 25228 5516 25280 5568
rect 10214 5414 10266 5466
rect 10278 5414 10330 5466
rect 10342 5414 10394 5466
rect 10406 5414 10458 5466
rect 10470 5414 10522 5466
rect 19478 5414 19530 5466
rect 19542 5414 19594 5466
rect 19606 5414 19658 5466
rect 19670 5414 19722 5466
rect 19734 5414 19786 5466
rect 9312 5355 9364 5364
rect 9312 5321 9321 5355
rect 9321 5321 9355 5355
rect 9355 5321 9364 5355
rect 9312 5312 9364 5321
rect 9680 5355 9732 5364
rect 9680 5321 9689 5355
rect 9689 5321 9723 5355
rect 9723 5321 9732 5355
rect 9680 5312 9732 5321
rect 8116 5244 8168 5296
rect 9864 5287 9916 5296
rect 9864 5253 9873 5287
rect 9873 5253 9907 5287
rect 9907 5253 9916 5287
rect 9864 5244 9916 5253
rect 9588 5219 9640 5228
rect 9588 5185 9597 5219
rect 9597 5185 9631 5219
rect 9631 5185 9640 5219
rect 9588 5176 9640 5185
rect 10140 5219 10192 5228
rect 10140 5185 10149 5219
rect 10149 5185 10183 5219
rect 10183 5185 10192 5219
rect 10140 5176 10192 5185
rect 11244 5312 11296 5364
rect 11520 5355 11572 5364
rect 11520 5321 11529 5355
rect 11529 5321 11563 5355
rect 11563 5321 11572 5355
rect 11520 5312 11572 5321
rect 11888 5312 11940 5364
rect 16120 5312 16172 5364
rect 12256 5244 12308 5296
rect 10692 5219 10744 5228
rect 10692 5185 10701 5219
rect 10701 5185 10735 5219
rect 10735 5185 10744 5219
rect 10692 5176 10744 5185
rect 10876 5176 10928 5228
rect 11796 5219 11848 5228
rect 11796 5185 11805 5219
rect 11805 5185 11839 5219
rect 11839 5185 11848 5219
rect 11796 5176 11848 5185
rect 10416 5151 10468 5160
rect 10416 5117 10425 5151
rect 10425 5117 10459 5151
rect 10459 5117 10468 5151
rect 10416 5108 10468 5117
rect 9956 5040 10008 5092
rect 12164 5176 12216 5228
rect 12900 5176 12952 5228
rect 13360 5176 13412 5228
rect 14004 5176 14056 5228
rect 14280 5176 14332 5228
rect 15292 5244 15344 5296
rect 12624 5151 12676 5160
rect 12624 5117 12633 5151
rect 12633 5117 12667 5151
rect 12667 5117 12676 5151
rect 12624 5108 12676 5117
rect 13084 5151 13136 5160
rect 13084 5117 13093 5151
rect 13093 5117 13127 5151
rect 13127 5117 13136 5151
rect 13084 5108 13136 5117
rect 13912 5151 13964 5160
rect 13912 5117 13921 5151
rect 13921 5117 13955 5151
rect 13955 5117 13964 5151
rect 13912 5108 13964 5117
rect 14556 5108 14608 5160
rect 17868 5312 17920 5364
rect 18328 5312 18380 5364
rect 19892 5312 19944 5364
rect 16764 5244 16816 5296
rect 17592 5244 17644 5296
rect 21640 5244 21692 5296
rect 16948 5219 17000 5228
rect 16948 5185 16982 5219
rect 16982 5185 17000 5219
rect 16948 5176 17000 5185
rect 18328 5219 18380 5228
rect 18328 5185 18337 5219
rect 18337 5185 18371 5219
rect 18371 5185 18380 5219
rect 18328 5176 18380 5185
rect 18604 5219 18656 5228
rect 18604 5185 18613 5219
rect 18613 5185 18647 5219
rect 18647 5185 18656 5219
rect 18604 5176 18656 5185
rect 19248 5176 19300 5228
rect 22008 5312 22060 5364
rect 22652 5287 22704 5296
rect 22652 5253 22661 5287
rect 22661 5253 22695 5287
rect 22695 5253 22704 5287
rect 22652 5244 22704 5253
rect 24032 5287 24084 5296
rect 24032 5253 24066 5287
rect 24066 5253 24084 5287
rect 24032 5244 24084 5253
rect 21916 5219 21968 5228
rect 21916 5185 21925 5219
rect 21925 5185 21959 5219
rect 21959 5185 21968 5219
rect 21916 5176 21968 5185
rect 21548 5108 21600 5160
rect 23020 5176 23072 5228
rect 24860 5176 24912 5228
rect 23572 5108 23624 5160
rect 10048 4972 10100 5024
rect 11060 4972 11112 5024
rect 11704 5015 11756 5024
rect 11704 4981 11713 5015
rect 11713 4981 11747 5015
rect 11747 4981 11756 5015
rect 11704 4972 11756 4981
rect 12440 4972 12492 5024
rect 12900 4972 12952 5024
rect 13176 5015 13228 5024
rect 13176 4981 13185 5015
rect 13185 4981 13219 5015
rect 13219 4981 13228 5015
rect 13176 4972 13228 4981
rect 13452 4972 13504 5024
rect 13544 4972 13596 5024
rect 14188 5015 14240 5024
rect 14188 4981 14197 5015
rect 14197 4981 14231 5015
rect 14231 4981 14240 5015
rect 14188 4972 14240 4981
rect 14740 5015 14792 5024
rect 14740 4981 14749 5015
rect 14749 4981 14783 5015
rect 14783 4981 14792 5015
rect 14740 4972 14792 4981
rect 15384 4972 15436 5024
rect 16120 4972 16172 5024
rect 17960 4972 18012 5024
rect 19248 4972 19300 5024
rect 23112 5015 23164 5024
rect 23112 4981 23121 5015
rect 23121 4981 23155 5015
rect 23155 4981 23164 5015
rect 23112 4972 23164 4981
rect 24492 4972 24544 5024
rect 25228 4972 25280 5024
rect 5582 4870 5634 4922
rect 5646 4870 5698 4922
rect 5710 4870 5762 4922
rect 5774 4870 5826 4922
rect 5838 4870 5890 4922
rect 14846 4870 14898 4922
rect 14910 4870 14962 4922
rect 14974 4870 15026 4922
rect 15038 4870 15090 4922
rect 15102 4870 15154 4922
rect 24110 4870 24162 4922
rect 24174 4870 24226 4922
rect 24238 4870 24290 4922
rect 24302 4870 24354 4922
rect 24366 4870 24418 4922
rect 10140 4768 10192 4820
rect 12624 4768 12676 4820
rect 12992 4768 13044 4820
rect 17408 4768 17460 4820
rect 18144 4811 18196 4820
rect 18144 4777 18153 4811
rect 18153 4777 18187 4811
rect 18187 4777 18196 4811
rect 18144 4768 18196 4777
rect 20536 4768 20588 4820
rect 23112 4768 23164 4820
rect 12256 4700 12308 4752
rect 13360 4700 13412 4752
rect 9312 4564 9364 4616
rect 10140 4632 10192 4684
rect 10416 4607 10468 4616
rect 10416 4573 10425 4607
rect 10425 4573 10459 4607
rect 10459 4573 10468 4607
rect 10416 4564 10468 4573
rect 11612 4632 11664 4684
rect 10784 4564 10836 4616
rect 11428 4607 11480 4616
rect 11428 4573 11437 4607
rect 11437 4573 11471 4607
rect 11471 4573 11480 4607
rect 11428 4564 11480 4573
rect 12164 4564 12216 4616
rect 12624 4564 12676 4616
rect 12900 4632 12952 4684
rect 14740 4632 14792 4684
rect 13176 4607 13228 4616
rect 13176 4573 13185 4607
rect 13185 4573 13219 4607
rect 13219 4573 13228 4607
rect 13176 4564 13228 4573
rect 14096 4607 14148 4616
rect 14096 4573 14105 4607
rect 14105 4573 14139 4607
rect 14139 4573 14148 4607
rect 14096 4564 14148 4573
rect 14556 4564 14608 4616
rect 16120 4607 16172 4616
rect 16120 4573 16129 4607
rect 16129 4573 16163 4607
rect 16163 4573 16172 4607
rect 16120 4564 16172 4573
rect 17224 4564 17276 4616
rect 18420 4607 18472 4616
rect 18420 4573 18429 4607
rect 18429 4573 18463 4607
rect 18463 4573 18472 4607
rect 18420 4564 18472 4573
rect 18972 4564 19024 4616
rect 21180 4632 21232 4684
rect 21916 4632 21968 4684
rect 23940 4700 23992 4752
rect 23020 4632 23072 4684
rect 15292 4496 15344 4548
rect 17776 4539 17828 4548
rect 17776 4505 17785 4539
rect 17785 4505 17819 4539
rect 17819 4505 17828 4539
rect 17776 4496 17828 4505
rect 18144 4496 18196 4548
rect 18788 4539 18840 4548
rect 18788 4505 18797 4539
rect 18797 4505 18831 4539
rect 18831 4505 18840 4539
rect 18788 4496 18840 4505
rect 20352 4564 20404 4616
rect 20536 4564 20588 4616
rect 21548 4607 21600 4616
rect 21548 4573 21557 4607
rect 21557 4573 21591 4607
rect 21591 4573 21600 4607
rect 21548 4564 21600 4573
rect 12624 4428 12676 4480
rect 16672 4471 16724 4480
rect 16672 4437 16681 4471
rect 16681 4437 16715 4471
rect 16715 4437 16724 4471
rect 16672 4428 16724 4437
rect 19340 4428 19392 4480
rect 19984 4496 20036 4548
rect 22560 4564 22612 4616
rect 22744 4607 22796 4616
rect 22744 4573 22753 4607
rect 22753 4573 22787 4607
rect 22787 4573 22796 4607
rect 22744 4564 22796 4573
rect 21824 4496 21876 4548
rect 22008 4496 22060 4548
rect 28356 4607 28408 4616
rect 28356 4573 28365 4607
rect 28365 4573 28399 4607
rect 28399 4573 28408 4607
rect 28356 4564 28408 4573
rect 20076 4428 20128 4480
rect 20628 4471 20680 4480
rect 20628 4437 20637 4471
rect 20637 4437 20671 4471
rect 20671 4437 20680 4471
rect 20628 4428 20680 4437
rect 10214 4326 10266 4378
rect 10278 4326 10330 4378
rect 10342 4326 10394 4378
rect 10406 4326 10458 4378
rect 10470 4326 10522 4378
rect 19478 4326 19530 4378
rect 19542 4326 19594 4378
rect 19606 4326 19658 4378
rect 19670 4326 19722 4378
rect 19734 4326 19786 4378
rect 8116 4088 8168 4140
rect 9956 4088 10008 4140
rect 11704 4224 11756 4276
rect 10600 4088 10652 4140
rect 12164 4088 12216 4140
rect 12256 4131 12308 4140
rect 12256 4097 12265 4131
rect 12265 4097 12299 4131
rect 12299 4097 12308 4131
rect 12808 4224 12860 4276
rect 14096 4224 14148 4276
rect 19340 4224 19392 4276
rect 21548 4224 21600 4276
rect 14188 4156 14240 4208
rect 17040 4156 17092 4208
rect 18972 4199 19024 4208
rect 12256 4088 12308 4097
rect 10784 4020 10836 4072
rect 12624 4131 12676 4140
rect 12624 4097 12633 4131
rect 12633 4097 12667 4131
rect 12667 4097 12676 4131
rect 12624 4088 12676 4097
rect 12900 4088 12952 4140
rect 13176 4088 13228 4140
rect 16672 4131 16724 4140
rect 16672 4097 16681 4131
rect 16681 4097 16715 4131
rect 16715 4097 16724 4131
rect 16672 4088 16724 4097
rect 17224 4131 17276 4140
rect 12992 4020 13044 4072
rect 15384 4063 15436 4072
rect 15384 4029 15393 4063
rect 15393 4029 15427 4063
rect 15427 4029 15436 4063
rect 15384 4020 15436 4029
rect 17224 4097 17233 4131
rect 17233 4097 17267 4131
rect 17267 4097 17276 4131
rect 17224 4088 17276 4097
rect 17408 4131 17460 4140
rect 17408 4097 17417 4131
rect 17417 4097 17451 4131
rect 17451 4097 17460 4131
rect 17408 4088 17460 4097
rect 17776 4088 17828 4140
rect 18972 4165 18981 4199
rect 18981 4165 19015 4199
rect 19015 4165 19024 4199
rect 18972 4156 19024 4165
rect 20628 4156 20680 4208
rect 21916 4156 21968 4208
rect 11428 3952 11480 4004
rect 10140 3884 10192 3936
rect 11612 3884 11664 3936
rect 11796 3884 11848 3936
rect 12164 3884 12216 3936
rect 12900 3884 12952 3936
rect 13268 3884 13320 3936
rect 16948 3927 17000 3936
rect 16948 3893 16957 3927
rect 16957 3893 16991 3927
rect 16991 3893 17000 3927
rect 16948 3884 17000 3893
rect 18144 4088 18196 4140
rect 19708 4088 19760 4140
rect 19892 4088 19944 4140
rect 18604 4020 18656 4072
rect 21916 4063 21968 4072
rect 21916 4029 21925 4063
rect 21925 4029 21959 4063
rect 21959 4029 21968 4063
rect 21916 4020 21968 4029
rect 23940 4131 23992 4140
rect 23940 4097 23958 4131
rect 23958 4097 23992 4131
rect 23940 4088 23992 4097
rect 22744 4020 22796 4072
rect 24492 4020 24544 4072
rect 19248 3884 19300 3936
rect 5582 3782 5634 3834
rect 5646 3782 5698 3834
rect 5710 3782 5762 3834
rect 5774 3782 5826 3834
rect 5838 3782 5890 3834
rect 14846 3782 14898 3834
rect 14910 3782 14962 3834
rect 14974 3782 15026 3834
rect 15038 3782 15090 3834
rect 15102 3782 15154 3834
rect 24110 3782 24162 3834
rect 24174 3782 24226 3834
rect 24238 3782 24290 3834
rect 24302 3782 24354 3834
rect 24366 3782 24418 3834
rect 13084 3680 13136 3732
rect 17776 3680 17828 3732
rect 18420 3680 18472 3732
rect 18972 3680 19024 3732
rect 12256 3612 12308 3664
rect 13268 3612 13320 3664
rect 13728 3655 13780 3664
rect 13728 3621 13737 3655
rect 13737 3621 13771 3655
rect 13771 3621 13780 3655
rect 13728 3612 13780 3621
rect 19248 3612 19300 3664
rect 21916 3680 21968 3732
rect 10876 3519 10928 3528
rect 10876 3485 10885 3519
rect 10885 3485 10919 3519
rect 10919 3485 10928 3519
rect 10876 3476 10928 3485
rect 11796 3476 11848 3528
rect 11888 3476 11940 3528
rect 12440 3544 12492 3596
rect 13176 3587 13228 3596
rect 11428 3451 11480 3460
rect 11428 3417 11437 3451
rect 11437 3417 11471 3451
rect 11471 3417 11480 3451
rect 11428 3408 11480 3417
rect 11612 3451 11664 3460
rect 11612 3417 11621 3451
rect 11621 3417 11655 3451
rect 11655 3417 11664 3451
rect 11612 3408 11664 3417
rect 10968 3383 11020 3392
rect 10968 3349 10983 3383
rect 10983 3349 11017 3383
rect 11017 3349 11020 3383
rect 10968 3340 11020 3349
rect 12624 3476 12676 3528
rect 13176 3553 13185 3587
rect 13185 3553 13219 3587
rect 13219 3553 13228 3587
rect 13176 3544 13228 3553
rect 13544 3544 13596 3596
rect 18604 3544 18656 3596
rect 13452 3519 13504 3528
rect 13452 3485 13461 3519
rect 13461 3485 13495 3519
rect 13495 3485 13504 3519
rect 13452 3476 13504 3485
rect 16764 3476 16816 3528
rect 17960 3476 18012 3528
rect 18144 3519 18196 3528
rect 18144 3485 18153 3519
rect 18153 3485 18187 3519
rect 18187 3485 18196 3519
rect 18144 3476 18196 3485
rect 19248 3519 19300 3528
rect 19248 3485 19257 3519
rect 19257 3485 19291 3519
rect 19291 3485 19300 3519
rect 19248 3476 19300 3485
rect 14004 3408 14056 3460
rect 16948 3408 17000 3460
rect 17408 3340 17460 3392
rect 19708 3519 19760 3528
rect 19708 3485 19717 3519
rect 19717 3485 19751 3519
rect 19751 3485 19760 3519
rect 19708 3476 19760 3485
rect 19892 3544 19944 3596
rect 21456 3476 21508 3528
rect 24492 3476 24544 3528
rect 20352 3408 20404 3460
rect 22836 3408 22888 3460
rect 19984 3340 20036 3392
rect 22284 3340 22336 3392
rect 28080 3340 28132 3392
rect 10214 3238 10266 3290
rect 10278 3238 10330 3290
rect 10342 3238 10394 3290
rect 10406 3238 10458 3290
rect 10470 3238 10522 3290
rect 19478 3238 19530 3290
rect 19542 3238 19594 3290
rect 19606 3238 19658 3290
rect 19670 3238 19722 3290
rect 19734 3238 19786 3290
rect 8208 3179 8260 3188
rect 8208 3145 8217 3179
rect 8217 3145 8251 3179
rect 8251 3145 8260 3179
rect 8208 3136 8260 3145
rect 11980 3136 12032 3188
rect 13176 3136 13228 3188
rect 20352 3179 20404 3188
rect 20352 3145 20361 3179
rect 20361 3145 20395 3179
rect 20395 3145 20404 3179
rect 20352 3136 20404 3145
rect 8116 3000 8168 3052
rect 10968 2932 11020 2984
rect 13728 3000 13780 3052
rect 15384 3068 15436 3120
rect 19892 3068 19944 3120
rect 20076 3000 20128 3052
rect 28080 3043 28132 3052
rect 28080 3009 28089 3043
rect 28089 3009 28123 3043
rect 28123 3009 28132 3043
rect 28080 3000 28132 3009
rect 13268 2864 13320 2916
rect 1676 2796 1728 2848
rect 5908 2796 5960 2848
rect 28264 2839 28316 2848
rect 28264 2805 28273 2839
rect 28273 2805 28307 2839
rect 28307 2805 28316 2839
rect 28264 2796 28316 2805
rect 5582 2694 5634 2746
rect 5646 2694 5698 2746
rect 5710 2694 5762 2746
rect 5774 2694 5826 2746
rect 5838 2694 5890 2746
rect 14846 2694 14898 2746
rect 14910 2694 14962 2746
rect 14974 2694 15026 2746
rect 15038 2694 15090 2746
rect 15102 2694 15154 2746
rect 24110 2694 24162 2746
rect 24174 2694 24226 2746
rect 24238 2694 24290 2746
rect 24302 2694 24354 2746
rect 24366 2694 24418 2746
rect 17040 2635 17092 2644
rect 17040 2601 17049 2635
rect 17049 2601 17083 2635
rect 17083 2601 17092 2635
rect 17040 2592 17092 2601
rect 20720 2635 20772 2644
rect 20720 2601 20729 2635
rect 20729 2601 20763 2635
rect 20763 2601 20772 2635
rect 20720 2592 20772 2601
rect 5908 2456 5960 2508
rect 20444 2524 20496 2576
rect 18512 2456 18564 2508
rect 20352 2456 20404 2508
rect 3240 2388 3292 2440
rect 6460 2388 6512 2440
rect 12256 2388 12308 2440
rect 1676 2363 1728 2372
rect 1676 2329 1685 2363
rect 1685 2329 1719 2363
rect 1719 2329 1728 2363
rect 1676 2320 1728 2329
rect 15660 2320 15712 2372
rect 16764 2320 16816 2372
rect 2228 2295 2280 2304
rect 2228 2261 2237 2295
rect 2237 2261 2271 2295
rect 2271 2261 2280 2295
rect 2228 2252 2280 2261
rect 5172 2252 5224 2304
rect 18696 2252 18748 2304
rect 20720 2388 20772 2440
rect 22284 2431 22336 2440
rect 22284 2397 22293 2431
rect 22293 2397 22327 2431
rect 22327 2397 22336 2431
rect 22284 2388 22336 2397
rect 25228 2431 25280 2440
rect 25228 2397 25237 2431
rect 25237 2397 25271 2431
rect 25271 2397 25280 2431
rect 25228 2388 25280 2397
rect 26424 2388 26476 2440
rect 21916 2252 21968 2304
rect 25136 2252 25188 2304
rect 27712 2252 27764 2304
rect 10214 2150 10266 2202
rect 10278 2150 10330 2202
rect 10342 2150 10394 2202
rect 10406 2150 10458 2202
rect 10470 2150 10522 2202
rect 19478 2150 19530 2202
rect 19542 2150 19594 2202
rect 19606 2150 19658 2202
rect 19670 2150 19722 2202
rect 19734 2150 19786 2202
<< metal2 >>
rect 662 29200 718 30000
rect 1306 29200 1362 30000
rect 2594 29322 2650 30000
rect 2424 29294 2650 29322
rect 1674 27976 1730 27985
rect 1674 27911 1730 27920
rect 1688 27470 1716 27911
rect 2424 27606 2452 29294
rect 2594 29200 2650 29294
rect 3882 29322 3938 30000
rect 3882 29294 4016 29322
rect 3882 29200 3938 29294
rect 3988 27606 4016 29294
rect 4526 29200 4582 30000
rect 5814 29200 5870 30000
rect 7102 29200 7158 30000
rect 8390 29200 8446 30000
rect 9034 29200 9090 30000
rect 10322 29322 10378 30000
rect 10322 29294 10548 29322
rect 10322 29200 10378 29294
rect 5582 27772 5890 27792
rect 5582 27770 5588 27772
rect 5644 27770 5668 27772
rect 5724 27770 5748 27772
rect 5804 27770 5828 27772
rect 5884 27770 5890 27772
rect 5644 27718 5646 27770
rect 5826 27718 5828 27770
rect 5582 27716 5588 27718
rect 5644 27716 5668 27718
rect 5724 27716 5748 27718
rect 5804 27716 5828 27718
rect 5884 27716 5890 27718
rect 5582 27696 5890 27716
rect 2412 27600 2464 27606
rect 2412 27542 2464 27548
rect 3976 27600 4028 27606
rect 3976 27542 4028 27548
rect 1676 27464 1728 27470
rect 1676 27406 1728 27412
rect 1688 27130 1716 27406
rect 3148 27396 3200 27402
rect 3148 27338 3200 27344
rect 1768 27328 1820 27334
rect 1768 27270 1820 27276
rect 1676 27124 1728 27130
rect 1676 27066 1728 27072
rect 1400 26988 1452 26994
rect 1400 26930 1452 26936
rect 1412 26625 1440 26930
rect 1584 26784 1636 26790
rect 1584 26726 1636 26732
rect 1398 26616 1454 26625
rect 1398 26551 1454 26560
rect 1400 26376 1452 26382
rect 1400 26318 1452 26324
rect 1412 25945 1440 26318
rect 1398 25936 1454 25945
rect 1398 25871 1454 25880
rect 1400 24812 1452 24818
rect 1400 24754 1452 24760
rect 1412 24585 1440 24754
rect 1398 24576 1454 24585
rect 1398 24511 1454 24520
rect 1400 23520 1452 23526
rect 1400 23462 1452 23468
rect 1412 23225 1440 23462
rect 1398 23216 1454 23225
rect 1398 23151 1454 23160
rect 1400 21344 1452 21350
rect 1400 21286 1452 21292
rect 1412 21185 1440 21286
rect 1398 21176 1454 21185
rect 1398 21111 1454 21120
rect 1400 19848 1452 19854
rect 1398 19816 1400 19825
rect 1452 19816 1454 19825
rect 1398 19751 1454 19760
rect 1412 19514 1440 19751
rect 1400 19508 1452 19514
rect 1400 19450 1452 19456
rect 1596 19174 1624 26726
rect 1676 24608 1728 24614
rect 1676 24550 1728 24556
rect 1584 19168 1636 19174
rect 1584 19110 1636 19116
rect 1400 18760 1452 18766
rect 1400 18702 1452 18708
rect 1412 18465 1440 18702
rect 1398 18456 1454 18465
rect 1398 18391 1454 18400
rect 1398 17096 1454 17105
rect 1398 17031 1400 17040
rect 1452 17031 1454 17040
rect 1400 17002 1452 17008
rect 1688 16574 1716 24550
rect 1780 17241 1808 27270
rect 3160 21078 3188 27338
rect 5582 26684 5890 26704
rect 5582 26682 5588 26684
rect 5644 26682 5668 26684
rect 5724 26682 5748 26684
rect 5804 26682 5828 26684
rect 5884 26682 5890 26684
rect 5644 26630 5646 26682
rect 5826 26630 5828 26682
rect 5582 26628 5588 26630
rect 5644 26628 5668 26630
rect 5724 26628 5748 26630
rect 5804 26628 5828 26630
rect 5884 26628 5890 26630
rect 5582 26608 5890 26628
rect 5582 25596 5890 25616
rect 5582 25594 5588 25596
rect 5644 25594 5668 25596
rect 5724 25594 5748 25596
rect 5804 25594 5828 25596
rect 5884 25594 5890 25596
rect 5644 25542 5646 25594
rect 5826 25542 5828 25594
rect 5582 25540 5588 25542
rect 5644 25540 5668 25542
rect 5724 25540 5748 25542
rect 5804 25540 5828 25542
rect 5884 25540 5890 25542
rect 5582 25520 5890 25540
rect 9048 24886 9076 29200
rect 10520 27470 10548 29294
rect 11610 29200 11666 30000
rect 12898 29200 12954 30000
rect 13542 29200 13598 30000
rect 14830 29200 14886 30000
rect 16118 29322 16174 30000
rect 16118 29294 16528 29322
rect 16118 29200 16174 29294
rect 14846 27772 15154 27792
rect 14846 27770 14852 27772
rect 14908 27770 14932 27772
rect 14988 27770 15012 27772
rect 15068 27770 15092 27772
rect 15148 27770 15154 27772
rect 14908 27718 14910 27770
rect 15090 27718 15092 27770
rect 14846 27716 14852 27718
rect 14908 27716 14932 27718
rect 14988 27716 15012 27718
rect 15068 27716 15092 27718
rect 15148 27716 15154 27718
rect 14846 27696 15154 27716
rect 16500 27606 16528 29294
rect 17406 29200 17462 30000
rect 18050 29200 18106 30000
rect 19338 29322 19394 30000
rect 19338 29294 19472 29322
rect 19338 29200 19394 29294
rect 19444 27606 19472 29294
rect 20626 29200 20682 30000
rect 21270 29200 21326 30000
rect 22558 29322 22614 30000
rect 22388 29294 22614 29322
rect 21284 27606 21312 29200
rect 22388 27606 22416 29294
rect 22558 29200 22614 29294
rect 23846 29322 23902 30000
rect 25134 29322 25190 30000
rect 25778 29322 25834 30000
rect 23846 29294 23980 29322
rect 23846 29200 23902 29294
rect 23952 27606 23980 29294
rect 25134 29294 25544 29322
rect 25134 29200 25190 29294
rect 24110 27772 24418 27792
rect 24110 27770 24116 27772
rect 24172 27770 24196 27772
rect 24252 27770 24276 27772
rect 24332 27770 24356 27772
rect 24412 27770 24418 27772
rect 24172 27718 24174 27770
rect 24354 27718 24356 27770
rect 24110 27716 24116 27718
rect 24172 27716 24196 27718
rect 24252 27716 24276 27718
rect 24332 27716 24356 27718
rect 24412 27716 24418 27718
rect 24110 27696 24418 27716
rect 25516 27606 25544 29294
rect 25778 29294 25912 29322
rect 25778 29200 25834 29294
rect 25884 27606 25912 29294
rect 27066 29200 27122 30000
rect 27526 29336 27582 29345
rect 28354 29322 28410 30000
rect 27526 29271 27582 29280
rect 28000 29294 28410 29322
rect 16488 27600 16540 27606
rect 16488 27542 16540 27548
rect 19432 27600 19484 27606
rect 19432 27542 19484 27548
rect 21272 27600 21324 27606
rect 21272 27542 21324 27548
rect 22376 27600 22428 27606
rect 22376 27542 22428 27548
rect 23940 27600 23992 27606
rect 23940 27542 23992 27548
rect 25504 27600 25556 27606
rect 25504 27542 25556 27548
rect 25872 27600 25924 27606
rect 25872 27542 25924 27548
rect 10508 27464 10560 27470
rect 10508 27406 10560 27412
rect 18328 27464 18380 27470
rect 18328 27406 18380 27412
rect 25136 27464 25188 27470
rect 25136 27406 25188 27412
rect 10784 27396 10836 27402
rect 10784 27338 10836 27344
rect 10214 27228 10522 27248
rect 10214 27226 10220 27228
rect 10276 27226 10300 27228
rect 10356 27226 10380 27228
rect 10436 27226 10460 27228
rect 10516 27226 10522 27228
rect 10276 27174 10278 27226
rect 10458 27174 10460 27226
rect 10214 27172 10220 27174
rect 10276 27172 10300 27174
rect 10356 27172 10380 27174
rect 10436 27172 10460 27174
rect 10516 27172 10522 27174
rect 10214 27152 10522 27172
rect 10214 26140 10522 26160
rect 10214 26138 10220 26140
rect 10276 26138 10300 26140
rect 10356 26138 10380 26140
rect 10436 26138 10460 26140
rect 10516 26138 10522 26140
rect 10276 26086 10278 26138
rect 10458 26086 10460 26138
rect 10214 26084 10220 26086
rect 10276 26084 10300 26086
rect 10356 26084 10380 26086
rect 10436 26084 10460 26086
rect 10516 26084 10522 26086
rect 10214 26064 10522 26084
rect 10214 25052 10522 25072
rect 10214 25050 10220 25052
rect 10276 25050 10300 25052
rect 10356 25050 10380 25052
rect 10436 25050 10460 25052
rect 10516 25050 10522 25052
rect 10276 24998 10278 25050
rect 10458 24998 10460 25050
rect 10214 24996 10220 24998
rect 10276 24996 10300 24998
rect 10356 24996 10380 24998
rect 10436 24996 10460 24998
rect 10516 24996 10522 24998
rect 10214 24976 10522 24996
rect 9036 24880 9088 24886
rect 9036 24822 9088 24828
rect 5582 24508 5890 24528
rect 5582 24506 5588 24508
rect 5644 24506 5668 24508
rect 5724 24506 5748 24508
rect 5804 24506 5828 24508
rect 5884 24506 5890 24508
rect 5644 24454 5646 24506
rect 5826 24454 5828 24506
rect 5582 24452 5588 24454
rect 5644 24452 5668 24454
rect 5724 24452 5748 24454
rect 5804 24452 5828 24454
rect 5884 24452 5890 24454
rect 5582 24432 5890 24452
rect 10214 23964 10522 23984
rect 10214 23962 10220 23964
rect 10276 23962 10300 23964
rect 10356 23962 10380 23964
rect 10436 23962 10460 23964
rect 10516 23962 10522 23964
rect 10276 23910 10278 23962
rect 10458 23910 10460 23962
rect 10214 23908 10220 23910
rect 10276 23908 10300 23910
rect 10356 23908 10380 23910
rect 10436 23908 10460 23910
rect 10516 23908 10522 23910
rect 10214 23888 10522 23908
rect 5582 23420 5890 23440
rect 5582 23418 5588 23420
rect 5644 23418 5668 23420
rect 5724 23418 5748 23420
rect 5804 23418 5828 23420
rect 5884 23418 5890 23420
rect 5644 23366 5646 23418
rect 5826 23366 5828 23418
rect 5582 23364 5588 23366
rect 5644 23364 5668 23366
rect 5724 23364 5748 23366
rect 5804 23364 5828 23366
rect 5884 23364 5890 23366
rect 5582 23344 5890 23364
rect 10214 22876 10522 22896
rect 10214 22874 10220 22876
rect 10276 22874 10300 22876
rect 10356 22874 10380 22876
rect 10436 22874 10460 22876
rect 10516 22874 10522 22876
rect 10276 22822 10278 22874
rect 10458 22822 10460 22874
rect 10214 22820 10220 22822
rect 10276 22820 10300 22822
rect 10356 22820 10380 22822
rect 10436 22820 10460 22822
rect 10516 22820 10522 22822
rect 10214 22800 10522 22820
rect 10508 22432 10560 22438
rect 10508 22374 10560 22380
rect 5582 22332 5890 22352
rect 5582 22330 5588 22332
rect 5644 22330 5668 22332
rect 5724 22330 5748 22332
rect 5804 22330 5828 22332
rect 5884 22330 5890 22332
rect 5644 22278 5646 22330
rect 5826 22278 5828 22330
rect 5582 22276 5588 22278
rect 5644 22276 5668 22278
rect 5724 22276 5748 22278
rect 5804 22276 5828 22278
rect 5884 22276 5890 22278
rect 5582 22256 5890 22276
rect 10520 22030 10548 22374
rect 7564 22024 7616 22030
rect 7564 21966 7616 21972
rect 9680 22024 9732 22030
rect 9680 21966 9732 21972
rect 10508 22024 10560 22030
rect 10508 21966 10560 21972
rect 6828 21548 6880 21554
rect 6828 21490 6880 21496
rect 5582 21244 5890 21264
rect 5582 21242 5588 21244
rect 5644 21242 5668 21244
rect 5724 21242 5748 21244
rect 5804 21242 5828 21244
rect 5884 21242 5890 21244
rect 5644 21190 5646 21242
rect 5826 21190 5828 21242
rect 5582 21188 5588 21190
rect 5644 21188 5668 21190
rect 5724 21188 5748 21190
rect 5804 21188 5828 21190
rect 5884 21188 5890 21190
rect 5582 21168 5890 21188
rect 3148 21072 3200 21078
rect 3148 21014 3200 21020
rect 6840 20398 6868 21490
rect 7576 21146 7604 21966
rect 7932 21888 7984 21894
rect 7932 21830 7984 21836
rect 9404 21888 9456 21894
rect 9404 21830 9456 21836
rect 7944 21554 7972 21830
rect 9416 21622 9444 21830
rect 9404 21616 9456 21622
rect 9404 21558 9456 21564
rect 7932 21548 7984 21554
rect 7932 21490 7984 21496
rect 9128 21480 9180 21486
rect 9128 21422 9180 21428
rect 7656 21344 7708 21350
rect 7656 21286 7708 21292
rect 9036 21344 9088 21350
rect 9036 21286 9088 21292
rect 7564 21140 7616 21146
rect 7564 21082 7616 21088
rect 7668 21078 7696 21286
rect 7656 21072 7708 21078
rect 7656 21014 7708 21020
rect 8116 21004 8168 21010
rect 8116 20946 8168 20952
rect 7104 20460 7156 20466
rect 7104 20402 7156 20408
rect 6828 20392 6880 20398
rect 6828 20334 6880 20340
rect 5582 20156 5890 20176
rect 5582 20154 5588 20156
rect 5644 20154 5668 20156
rect 5724 20154 5748 20156
rect 5804 20154 5828 20156
rect 5884 20154 5890 20156
rect 5644 20102 5646 20154
rect 5826 20102 5828 20154
rect 5582 20100 5588 20102
rect 5644 20100 5668 20102
rect 5724 20100 5748 20102
rect 5804 20100 5828 20102
rect 5884 20100 5890 20102
rect 5582 20080 5890 20100
rect 7116 20058 7144 20402
rect 7104 20052 7156 20058
rect 7104 19994 7156 20000
rect 8128 19922 8156 20946
rect 8208 20936 8260 20942
rect 8208 20878 8260 20884
rect 8220 20262 8248 20878
rect 9048 20874 9076 21286
rect 9036 20868 9088 20874
rect 9036 20810 9088 20816
rect 9140 20262 9168 21422
rect 9404 21072 9456 21078
rect 9404 21014 9456 21020
rect 9416 20398 9444 21014
rect 9496 20800 9548 20806
rect 9496 20742 9548 20748
rect 9508 20466 9536 20742
rect 9692 20602 9720 21966
rect 10140 21956 10192 21962
rect 10140 21898 10192 21904
rect 9772 21684 9824 21690
rect 9772 21626 9824 21632
rect 9784 20942 9812 21626
rect 9772 20936 9824 20942
rect 9772 20878 9824 20884
rect 9680 20596 9732 20602
rect 9680 20538 9732 20544
rect 10152 20534 10180 21898
rect 10520 21876 10548 21966
rect 10520 21848 10640 21876
rect 10214 21788 10522 21808
rect 10214 21786 10220 21788
rect 10276 21786 10300 21788
rect 10356 21786 10380 21788
rect 10436 21786 10460 21788
rect 10516 21786 10522 21788
rect 10276 21734 10278 21786
rect 10458 21734 10460 21786
rect 10214 21732 10220 21734
rect 10276 21732 10300 21734
rect 10356 21732 10380 21734
rect 10436 21732 10460 21734
rect 10516 21732 10522 21734
rect 10214 21712 10522 21732
rect 10214 20700 10522 20720
rect 10214 20698 10220 20700
rect 10276 20698 10300 20700
rect 10356 20698 10380 20700
rect 10436 20698 10460 20700
rect 10516 20698 10522 20700
rect 10276 20646 10278 20698
rect 10458 20646 10460 20698
rect 10214 20644 10220 20646
rect 10276 20644 10300 20646
rect 10356 20644 10380 20646
rect 10436 20644 10460 20646
rect 10516 20644 10522 20646
rect 10214 20624 10522 20644
rect 10140 20528 10192 20534
rect 10140 20470 10192 20476
rect 9496 20460 9548 20466
rect 9496 20402 9548 20408
rect 10048 20460 10100 20466
rect 10048 20402 10100 20408
rect 9404 20392 9456 20398
rect 9404 20334 9456 20340
rect 8208 20256 8260 20262
rect 8208 20198 8260 20204
rect 9128 20256 9180 20262
rect 9128 20198 9180 20204
rect 8116 19916 8168 19922
rect 8116 19858 8168 19864
rect 7748 19780 7800 19786
rect 7748 19722 7800 19728
rect 6920 19508 6972 19514
rect 6920 19450 6972 19456
rect 5582 19068 5890 19088
rect 5582 19066 5588 19068
rect 5644 19066 5668 19068
rect 5724 19066 5748 19068
rect 5804 19066 5828 19068
rect 5884 19066 5890 19068
rect 5644 19014 5646 19066
rect 5826 19014 5828 19066
rect 5582 19012 5588 19014
rect 5644 19012 5668 19014
rect 5724 19012 5748 19014
rect 5804 19012 5828 19014
rect 5884 19012 5890 19014
rect 5582 18992 5890 19012
rect 6932 18766 6960 19450
rect 7012 19372 7064 19378
rect 7012 19314 7064 19320
rect 6644 18760 6696 18766
rect 6644 18702 6696 18708
rect 6920 18760 6972 18766
rect 6920 18702 6972 18708
rect 6000 18216 6052 18222
rect 6000 18158 6052 18164
rect 4620 18080 4672 18086
rect 4620 18022 4672 18028
rect 1766 17232 1822 17241
rect 1766 17167 1822 17176
rect 4632 16590 4660 18022
rect 5582 17980 5890 18000
rect 5582 17978 5588 17980
rect 5644 17978 5668 17980
rect 5724 17978 5748 17980
rect 5804 17978 5828 17980
rect 5884 17978 5890 17980
rect 5644 17926 5646 17978
rect 5826 17926 5828 17978
rect 5582 17924 5588 17926
rect 5644 17924 5668 17926
rect 5724 17924 5748 17926
rect 5804 17924 5828 17926
rect 5884 17924 5890 17926
rect 5582 17904 5890 17924
rect 6012 17678 6040 18158
rect 6656 18154 6684 18702
rect 7024 18426 7052 19314
rect 7288 18760 7340 18766
rect 7288 18702 7340 18708
rect 7012 18420 7064 18426
rect 7012 18362 7064 18368
rect 7300 18222 7328 18702
rect 6736 18216 6788 18222
rect 6736 18158 6788 18164
rect 7288 18216 7340 18222
rect 7288 18158 7340 18164
rect 7380 18216 7432 18222
rect 7380 18158 7432 18164
rect 6644 18148 6696 18154
rect 6644 18090 6696 18096
rect 6748 18086 6776 18158
rect 6736 18080 6788 18086
rect 6736 18022 6788 18028
rect 6000 17672 6052 17678
rect 6000 17614 6052 17620
rect 5582 16892 5890 16912
rect 5582 16890 5588 16892
rect 5644 16890 5668 16892
rect 5724 16890 5748 16892
rect 5804 16890 5828 16892
rect 5884 16890 5890 16892
rect 5644 16838 5646 16890
rect 5826 16838 5828 16890
rect 5582 16836 5588 16838
rect 5644 16836 5668 16838
rect 5724 16836 5748 16838
rect 5804 16836 5828 16838
rect 5884 16836 5890 16838
rect 5582 16816 5890 16836
rect 4620 16584 4672 16590
rect 1688 16546 1808 16574
rect 1492 16448 1544 16454
rect 1490 16416 1492 16425
rect 1544 16416 1546 16425
rect 1490 16351 1546 16360
rect 1400 13864 1452 13870
rect 1400 13806 1452 13812
rect 1412 13705 1440 13806
rect 1398 13696 1454 13705
rect 1398 13631 1454 13640
rect 1400 10464 1452 10470
rect 1400 10406 1452 10412
rect 1412 10305 1440 10406
rect 1398 10296 1454 10305
rect 1398 10231 1454 10240
rect 1674 8936 1730 8945
rect 1674 8871 1676 8880
rect 1728 8871 1730 8880
rect 1676 8842 1728 8848
rect 1400 8492 1452 8498
rect 1400 8434 1452 8440
rect 1412 8265 1440 8434
rect 1780 8401 1808 16546
rect 4620 16526 4672 16532
rect 5908 16108 5960 16114
rect 5908 16050 5960 16056
rect 5172 15904 5224 15910
rect 5172 15846 5224 15852
rect 5184 15502 5212 15846
rect 5582 15804 5890 15824
rect 5582 15802 5588 15804
rect 5644 15802 5668 15804
rect 5724 15802 5748 15804
rect 5804 15802 5828 15804
rect 5884 15802 5890 15804
rect 5644 15750 5646 15802
rect 5826 15750 5828 15802
rect 5582 15748 5588 15750
rect 5644 15748 5668 15750
rect 5724 15748 5748 15750
rect 5804 15748 5828 15750
rect 5884 15748 5890 15750
rect 5582 15728 5890 15748
rect 5920 15706 5948 16050
rect 5908 15700 5960 15706
rect 5908 15642 5960 15648
rect 5172 15496 5224 15502
rect 5172 15438 5224 15444
rect 5632 15496 5684 15502
rect 5632 15438 5684 15444
rect 5644 15026 5672 15438
rect 6012 15026 6040 17614
rect 6092 17604 6144 17610
rect 6092 17546 6144 17552
rect 6104 17338 6132 17546
rect 6748 17490 6776 18022
rect 7392 17542 7420 18158
rect 6656 17462 6776 17490
rect 7380 17536 7432 17542
rect 7380 17478 7432 17484
rect 6092 17332 6144 17338
rect 6092 17274 6144 17280
rect 6656 17134 6684 17462
rect 7392 17270 7420 17478
rect 7380 17264 7432 17270
rect 7380 17206 7432 17212
rect 6644 17128 6696 17134
rect 6644 17070 6696 17076
rect 7472 17128 7524 17134
rect 7472 17070 7524 17076
rect 6656 16114 6684 17070
rect 7484 16794 7512 17070
rect 7472 16788 7524 16794
rect 7472 16730 7524 16736
rect 7656 16788 7708 16794
rect 7656 16730 7708 16736
rect 7668 16250 7696 16730
rect 7656 16244 7708 16250
rect 7656 16186 7708 16192
rect 6644 16108 6696 16114
rect 6644 16050 6696 16056
rect 7656 15972 7708 15978
rect 7656 15914 7708 15920
rect 7668 15638 7696 15914
rect 7656 15632 7708 15638
rect 7656 15574 7708 15580
rect 7288 15564 7340 15570
rect 7288 15506 7340 15512
rect 7196 15428 7248 15434
rect 7196 15370 7248 15376
rect 5632 15020 5684 15026
rect 5632 14962 5684 14968
rect 6000 15020 6052 15026
rect 6000 14962 6052 14968
rect 5582 14716 5890 14736
rect 5582 14714 5588 14716
rect 5644 14714 5668 14716
rect 5724 14714 5748 14716
rect 5804 14714 5828 14716
rect 5884 14714 5890 14716
rect 5644 14662 5646 14714
rect 5826 14662 5828 14714
rect 5582 14660 5588 14662
rect 5644 14660 5668 14662
rect 5724 14660 5748 14662
rect 5804 14660 5828 14662
rect 5884 14660 5890 14662
rect 5582 14640 5890 14660
rect 4436 14408 4488 14414
rect 4436 14350 4488 14356
rect 4448 13870 4476 14350
rect 6920 14340 6972 14346
rect 6920 14282 6972 14288
rect 6932 14074 6960 14282
rect 6920 14068 6972 14074
rect 6920 14010 6972 14016
rect 6552 14000 6604 14006
rect 6552 13942 6604 13948
rect 6276 13932 6328 13938
rect 6276 13874 6328 13880
rect 4436 13864 4488 13870
rect 4436 13806 4488 13812
rect 4448 12850 4476 13806
rect 5582 13628 5890 13648
rect 5582 13626 5588 13628
rect 5644 13626 5668 13628
rect 5724 13626 5748 13628
rect 5804 13626 5828 13628
rect 5884 13626 5890 13628
rect 5644 13574 5646 13626
rect 5826 13574 5828 13626
rect 5582 13572 5588 13574
rect 5644 13572 5668 13574
rect 5724 13572 5748 13574
rect 5804 13572 5828 13574
rect 5884 13572 5890 13574
rect 5582 13552 5890 13572
rect 6288 13530 6316 13874
rect 6564 13530 6592 13942
rect 7104 13932 7156 13938
rect 7104 13874 7156 13880
rect 6736 13864 6788 13870
rect 6736 13806 6788 13812
rect 6276 13524 6328 13530
rect 6276 13466 6328 13472
rect 6552 13524 6604 13530
rect 6552 13466 6604 13472
rect 6748 13326 6776 13806
rect 7012 13728 7064 13734
rect 7012 13670 7064 13676
rect 6828 13388 6880 13394
rect 6828 13330 6880 13336
rect 6736 13320 6788 13326
rect 6736 13262 6788 13268
rect 6736 12980 6788 12986
rect 6736 12922 6788 12928
rect 4436 12844 4488 12850
rect 4436 12786 4488 12792
rect 5908 12844 5960 12850
rect 5908 12786 5960 12792
rect 5582 12540 5890 12560
rect 5582 12538 5588 12540
rect 5644 12538 5668 12540
rect 5724 12538 5748 12540
rect 5804 12538 5828 12540
rect 5884 12538 5890 12540
rect 5644 12486 5646 12538
rect 5826 12486 5828 12538
rect 5582 12484 5588 12486
rect 5644 12484 5668 12486
rect 5724 12484 5748 12486
rect 5804 12484 5828 12486
rect 5884 12484 5890 12486
rect 5582 12464 5890 12484
rect 5920 12442 5948 12786
rect 6092 12640 6144 12646
rect 6092 12582 6144 12588
rect 5908 12436 5960 12442
rect 5908 12378 5960 12384
rect 6000 12232 6052 12238
rect 6000 12174 6052 12180
rect 6012 11762 6040 12174
rect 6104 12170 6132 12582
rect 6644 12368 6696 12374
rect 6644 12310 6696 12316
rect 6656 12238 6684 12310
rect 6644 12232 6696 12238
rect 6644 12174 6696 12180
rect 6092 12164 6144 12170
rect 6092 12106 6144 12112
rect 6552 12164 6604 12170
rect 6552 12106 6604 12112
rect 4528 11756 4580 11762
rect 4528 11698 4580 11704
rect 6000 11756 6052 11762
rect 6000 11698 6052 11704
rect 4540 11354 4568 11698
rect 5448 11552 5500 11558
rect 5448 11494 5500 11500
rect 4528 11348 4580 11354
rect 4528 11290 4580 11296
rect 5460 11234 5488 11494
rect 5582 11452 5890 11472
rect 5582 11450 5588 11452
rect 5644 11450 5668 11452
rect 5724 11450 5748 11452
rect 5804 11450 5828 11452
rect 5884 11450 5890 11452
rect 5644 11398 5646 11450
rect 5826 11398 5828 11450
rect 5582 11396 5588 11398
rect 5644 11396 5668 11398
rect 5724 11396 5748 11398
rect 5804 11396 5828 11398
rect 5884 11396 5890 11398
rect 5582 11376 5890 11396
rect 6564 11354 6592 12106
rect 6552 11348 6604 11354
rect 6552 11290 6604 11296
rect 5460 11206 5580 11234
rect 5552 11082 5580 11206
rect 5908 11144 5960 11150
rect 5908 11086 5960 11092
rect 5540 11076 5592 11082
rect 5540 11018 5592 11024
rect 5448 10464 5500 10470
rect 5448 10406 5500 10412
rect 5460 9994 5488 10406
rect 5582 10364 5890 10384
rect 5582 10362 5588 10364
rect 5644 10362 5668 10364
rect 5724 10362 5748 10364
rect 5804 10362 5828 10364
rect 5884 10362 5890 10364
rect 5644 10310 5646 10362
rect 5826 10310 5828 10362
rect 5582 10308 5588 10310
rect 5644 10308 5668 10310
rect 5724 10308 5748 10310
rect 5804 10308 5828 10310
rect 5884 10308 5890 10310
rect 5582 10288 5890 10308
rect 5920 10062 5948 11086
rect 6656 10826 6684 12174
rect 6748 12170 6776 12922
rect 6840 12646 6868 13330
rect 7024 12866 7052 13670
rect 7116 13530 7144 13874
rect 7104 13524 7156 13530
rect 7104 13466 7156 13472
rect 7104 12912 7156 12918
rect 6932 12860 7104 12866
rect 6932 12854 7156 12860
rect 6932 12838 7144 12854
rect 6828 12640 6880 12646
rect 6828 12582 6880 12588
rect 6840 12306 6868 12582
rect 6932 12442 6960 12838
rect 7012 12640 7064 12646
rect 7012 12582 7064 12588
rect 7024 12442 7052 12582
rect 6920 12436 6972 12442
rect 6920 12378 6972 12384
rect 7012 12436 7064 12442
rect 7012 12378 7064 12384
rect 6828 12300 6880 12306
rect 6828 12242 6880 12248
rect 6736 12164 6788 12170
rect 6736 12106 6788 12112
rect 7012 12096 7064 12102
rect 7012 12038 7064 12044
rect 7024 11694 7052 12038
rect 7104 11892 7156 11898
rect 7104 11834 7156 11840
rect 7012 11688 7064 11694
rect 7012 11630 7064 11636
rect 6828 11552 6880 11558
rect 6828 11494 6880 11500
rect 6840 11082 6868 11494
rect 7024 11354 7052 11630
rect 7012 11348 7064 11354
rect 7012 11290 7064 11296
rect 7116 11150 7144 11834
rect 7208 11218 7236 15370
rect 7196 11212 7248 11218
rect 7196 11154 7248 11160
rect 7104 11144 7156 11150
rect 7104 11086 7156 11092
rect 6828 11076 6880 11082
rect 6828 11018 6880 11024
rect 6656 10798 6960 10826
rect 6000 10668 6052 10674
rect 6000 10610 6052 10616
rect 5908 10056 5960 10062
rect 5908 9998 5960 10004
rect 5448 9988 5500 9994
rect 5448 9930 5500 9936
rect 6012 9382 6040 10610
rect 6932 10538 6960 10798
rect 7208 10742 7236 11154
rect 7196 10736 7248 10742
rect 7196 10678 7248 10684
rect 7104 10668 7156 10674
rect 7104 10610 7156 10616
rect 6920 10532 6972 10538
rect 6920 10474 6972 10480
rect 6828 10464 6880 10470
rect 6828 10406 6880 10412
rect 6840 10198 6868 10406
rect 6828 10192 6880 10198
rect 6828 10134 6880 10140
rect 6932 9450 6960 10474
rect 7116 10470 7144 10610
rect 7104 10464 7156 10470
rect 7104 10406 7156 10412
rect 7300 10266 7328 15506
rect 7668 15502 7696 15574
rect 7760 15502 7788 19722
rect 8128 18834 8156 19858
rect 8220 19718 8248 20198
rect 9140 19854 9168 20198
rect 8300 19848 8352 19854
rect 8300 19790 8352 19796
rect 9036 19848 9088 19854
rect 9036 19790 9088 19796
rect 9128 19848 9180 19854
rect 9128 19790 9180 19796
rect 8208 19712 8260 19718
rect 8208 19654 8260 19660
rect 8220 19446 8248 19654
rect 8208 19440 8260 19446
rect 8208 19382 8260 19388
rect 8312 19310 8340 19790
rect 8852 19372 8904 19378
rect 8852 19314 8904 19320
rect 8300 19304 8352 19310
rect 8300 19246 8352 19252
rect 8864 18970 8892 19314
rect 8852 18964 8904 18970
rect 8852 18906 8904 18912
rect 8116 18828 8168 18834
rect 8116 18770 8168 18776
rect 7840 18624 7892 18630
rect 7840 18566 7892 18572
rect 7852 18426 7880 18566
rect 7840 18420 7892 18426
rect 7840 18362 7892 18368
rect 8128 18222 8156 18770
rect 9048 18426 9076 19790
rect 9312 19780 9364 19786
rect 9312 19722 9364 19728
rect 9324 19514 9352 19722
rect 9312 19508 9364 19514
rect 9312 19450 9364 19456
rect 9416 19310 9444 20334
rect 9680 19712 9732 19718
rect 9680 19654 9732 19660
rect 9404 19304 9456 19310
rect 9404 19246 9456 19252
rect 9692 18766 9720 19654
rect 10060 19514 10088 20402
rect 10214 19612 10522 19632
rect 10214 19610 10220 19612
rect 10276 19610 10300 19612
rect 10356 19610 10380 19612
rect 10436 19610 10460 19612
rect 10516 19610 10522 19612
rect 10276 19558 10278 19610
rect 10458 19558 10460 19610
rect 10214 19556 10220 19558
rect 10276 19556 10300 19558
rect 10356 19556 10380 19558
rect 10436 19556 10460 19558
rect 10516 19556 10522 19558
rect 10214 19536 10522 19556
rect 10048 19508 10100 19514
rect 10048 19450 10100 19456
rect 9680 18760 9732 18766
rect 9680 18702 9732 18708
rect 9588 18692 9640 18698
rect 9588 18634 9640 18640
rect 9600 18426 9628 18634
rect 10214 18524 10522 18544
rect 10214 18522 10220 18524
rect 10276 18522 10300 18524
rect 10356 18522 10380 18524
rect 10436 18522 10460 18524
rect 10516 18522 10522 18524
rect 10276 18470 10278 18522
rect 10458 18470 10460 18522
rect 10214 18468 10220 18470
rect 10276 18468 10300 18470
rect 10356 18468 10380 18470
rect 10436 18468 10460 18470
rect 10516 18468 10522 18470
rect 10214 18448 10522 18468
rect 9036 18420 9088 18426
rect 9036 18362 9088 18368
rect 9588 18420 9640 18426
rect 9588 18362 9640 18368
rect 9680 18420 9732 18426
rect 9680 18362 9732 18368
rect 8116 18216 8168 18222
rect 8116 18158 8168 18164
rect 8128 17882 8156 18158
rect 8116 17876 8168 17882
rect 8116 17818 8168 17824
rect 9048 17678 9076 18362
rect 9692 18222 9720 18362
rect 9864 18352 9916 18358
rect 9864 18294 9916 18300
rect 9680 18216 9732 18222
rect 9680 18158 9732 18164
rect 9772 18216 9824 18222
rect 9772 18158 9824 18164
rect 9128 18080 9180 18086
rect 9128 18022 9180 18028
rect 9036 17672 9088 17678
rect 9036 17614 9088 17620
rect 8024 17604 8076 17610
rect 8024 17546 8076 17552
rect 8668 17604 8720 17610
rect 8668 17546 8720 17552
rect 8036 17134 8064 17546
rect 8680 17338 8708 17546
rect 8668 17332 8720 17338
rect 8668 17274 8720 17280
rect 7840 17128 7892 17134
rect 7840 17070 7892 17076
rect 8024 17128 8076 17134
rect 8024 17070 8076 17076
rect 7852 16046 7880 17070
rect 9048 16658 9076 17614
rect 9140 17202 9168 18022
rect 9128 17196 9180 17202
rect 9128 17138 9180 17144
rect 9312 17128 9364 17134
rect 9312 17070 9364 17076
rect 9036 16652 9088 16658
rect 9036 16594 9088 16600
rect 9324 16590 9352 17070
rect 9784 16590 9812 18158
rect 9876 17338 9904 18294
rect 10324 18284 10376 18290
rect 10324 18226 10376 18232
rect 10336 17814 10364 18226
rect 10612 17882 10640 21848
rect 10692 18624 10744 18630
rect 10692 18566 10744 18572
rect 10704 18290 10732 18566
rect 10692 18284 10744 18290
rect 10692 18226 10744 18232
rect 10600 17876 10652 17882
rect 10600 17818 10652 17824
rect 10324 17808 10376 17814
rect 10324 17750 10376 17756
rect 10214 17436 10522 17456
rect 10214 17434 10220 17436
rect 10276 17434 10300 17436
rect 10356 17434 10380 17436
rect 10436 17434 10460 17436
rect 10516 17434 10522 17436
rect 10276 17382 10278 17434
rect 10458 17382 10460 17434
rect 10214 17380 10220 17382
rect 10276 17380 10300 17382
rect 10356 17380 10380 17382
rect 10436 17380 10460 17382
rect 10516 17380 10522 17382
rect 10214 17360 10522 17380
rect 9864 17332 9916 17338
rect 9864 17274 9916 17280
rect 9876 16794 9904 17274
rect 10612 17270 10640 17818
rect 10600 17264 10652 17270
rect 10600 17206 10652 17212
rect 10324 16992 10376 16998
rect 10796 16946 10824 27338
rect 14846 26684 15154 26704
rect 14846 26682 14852 26684
rect 14908 26682 14932 26684
rect 14988 26682 15012 26684
rect 15068 26682 15092 26684
rect 15148 26682 15154 26684
rect 14908 26630 14910 26682
rect 15090 26630 15092 26682
rect 14846 26628 14852 26630
rect 14908 26628 14932 26630
rect 14988 26628 15012 26630
rect 15068 26628 15092 26630
rect 15148 26628 15154 26630
rect 14846 26608 15154 26628
rect 14846 25596 15154 25616
rect 14846 25594 14852 25596
rect 14908 25594 14932 25596
rect 14988 25594 15012 25596
rect 15068 25594 15092 25596
rect 15148 25594 15154 25596
rect 14908 25542 14910 25594
rect 15090 25542 15092 25594
rect 14846 25540 14852 25542
rect 14908 25540 14932 25542
rect 14988 25540 15012 25542
rect 15068 25540 15092 25542
rect 15148 25540 15154 25542
rect 14846 25520 15154 25540
rect 12164 24880 12216 24886
rect 12164 24822 12216 24828
rect 10876 22636 10928 22642
rect 10876 22578 10928 22584
rect 10888 20942 10916 22578
rect 11612 21956 11664 21962
rect 11612 21898 11664 21904
rect 11152 21548 11204 21554
rect 11152 21490 11204 21496
rect 10876 20936 10928 20942
rect 10876 20878 10928 20884
rect 10888 20466 10916 20878
rect 11164 20602 11192 21490
rect 11336 21344 11388 21350
rect 11336 21286 11388 21292
rect 11520 21344 11572 21350
rect 11520 21286 11572 21292
rect 11348 20874 11376 21286
rect 11532 21010 11560 21286
rect 11624 21146 11652 21898
rect 11612 21140 11664 21146
rect 11612 21082 11664 21088
rect 11520 21004 11572 21010
rect 11520 20946 11572 20952
rect 11244 20868 11296 20874
rect 11244 20810 11296 20816
rect 11336 20868 11388 20874
rect 11336 20810 11388 20816
rect 11256 20602 11284 20810
rect 11152 20596 11204 20602
rect 11152 20538 11204 20544
rect 11244 20596 11296 20602
rect 11244 20538 11296 20544
rect 10876 20460 10928 20466
rect 10876 20402 10928 20408
rect 11704 20256 11756 20262
rect 11704 20198 11756 20204
rect 11520 19780 11572 19786
rect 11520 19722 11572 19728
rect 11532 19514 11560 19722
rect 11520 19508 11572 19514
rect 11520 19450 11572 19456
rect 11716 19378 11744 20198
rect 11704 19372 11756 19378
rect 11704 19314 11756 19320
rect 10968 19304 11020 19310
rect 10968 19246 11020 19252
rect 11244 19304 11296 19310
rect 11244 19246 11296 19252
rect 10876 18964 10928 18970
rect 10876 18906 10928 18912
rect 10324 16934 10376 16940
rect 9864 16788 9916 16794
rect 9864 16730 9916 16736
rect 10336 16658 10364 16934
rect 10612 16918 10824 16946
rect 10324 16652 10376 16658
rect 10324 16594 10376 16600
rect 9312 16584 9364 16590
rect 9312 16526 9364 16532
rect 9772 16584 9824 16590
rect 9772 16526 9824 16532
rect 8300 16516 8352 16522
rect 8300 16458 8352 16464
rect 7840 16040 7892 16046
rect 7840 15982 7892 15988
rect 7852 15570 7880 15982
rect 8312 15706 8340 16458
rect 9220 16448 9272 16454
rect 9220 16390 9272 16396
rect 9232 16114 9260 16390
rect 9312 16244 9364 16250
rect 9312 16186 9364 16192
rect 9220 16108 9272 16114
rect 9220 16050 9272 16056
rect 9324 16046 9352 16186
rect 9784 16182 9812 16526
rect 10214 16348 10522 16368
rect 10214 16346 10220 16348
rect 10276 16346 10300 16348
rect 10356 16346 10380 16348
rect 10436 16346 10460 16348
rect 10516 16346 10522 16348
rect 10276 16294 10278 16346
rect 10458 16294 10460 16346
rect 10214 16292 10220 16294
rect 10276 16292 10300 16294
rect 10356 16292 10380 16294
rect 10436 16292 10460 16294
rect 10516 16292 10522 16294
rect 10214 16272 10522 16292
rect 9772 16176 9824 16182
rect 9772 16118 9824 16124
rect 9588 16108 9640 16114
rect 9588 16050 9640 16056
rect 9312 16040 9364 16046
rect 9312 15982 9364 15988
rect 8484 15904 8536 15910
rect 8484 15846 8536 15852
rect 9036 15904 9088 15910
rect 9036 15846 9088 15852
rect 8300 15700 8352 15706
rect 8300 15642 8352 15648
rect 7840 15564 7892 15570
rect 7840 15506 7892 15512
rect 8496 15502 8524 15846
rect 9048 15502 9076 15846
rect 7656 15496 7708 15502
rect 7656 15438 7708 15444
rect 7748 15496 7800 15502
rect 7748 15438 7800 15444
rect 8484 15496 8536 15502
rect 8484 15438 8536 15444
rect 9036 15496 9088 15502
rect 9036 15438 9088 15444
rect 8208 15088 8260 15094
rect 8208 15030 8260 15036
rect 8116 15020 8168 15026
rect 8116 14962 8168 14968
rect 8128 14074 8156 14962
rect 8116 14068 8168 14074
rect 8116 14010 8168 14016
rect 8024 14000 8076 14006
rect 8024 13942 8076 13948
rect 7932 13524 7984 13530
rect 7932 13466 7984 13472
rect 7656 13456 7708 13462
rect 7656 13398 7708 13404
rect 7380 13320 7432 13326
rect 7380 13262 7432 13268
rect 7392 12374 7420 13262
rect 7472 13184 7524 13190
rect 7472 13126 7524 13132
rect 7484 12986 7512 13126
rect 7472 12980 7524 12986
rect 7472 12922 7524 12928
rect 7472 12844 7524 12850
rect 7472 12786 7524 12792
rect 7380 12368 7432 12374
rect 7380 12310 7432 12316
rect 7484 12170 7512 12786
rect 7564 12232 7616 12238
rect 7564 12174 7616 12180
rect 7472 12164 7524 12170
rect 7472 12106 7524 12112
rect 7484 11830 7512 12106
rect 7472 11824 7524 11830
rect 7472 11766 7524 11772
rect 7380 11756 7432 11762
rect 7380 11698 7432 11704
rect 7392 11642 7420 11698
rect 7576 11694 7604 12174
rect 7668 11762 7696 13398
rect 7944 12986 7972 13466
rect 7932 12980 7984 12986
rect 7932 12922 7984 12928
rect 8036 12782 8064 13942
rect 8116 13864 8168 13870
rect 8116 13806 8168 13812
rect 8128 13530 8156 13806
rect 8220 13734 8248 15030
rect 9324 15026 9352 15982
rect 9600 15706 9628 16050
rect 9588 15700 9640 15706
rect 9588 15642 9640 15648
rect 10214 15260 10522 15280
rect 10214 15258 10220 15260
rect 10276 15258 10300 15260
rect 10356 15258 10380 15260
rect 10436 15258 10460 15260
rect 10516 15258 10522 15260
rect 10276 15206 10278 15258
rect 10458 15206 10460 15258
rect 10214 15204 10220 15206
rect 10276 15204 10300 15206
rect 10356 15204 10380 15206
rect 10436 15204 10460 15206
rect 10516 15204 10522 15206
rect 10214 15184 10522 15204
rect 10612 15094 10640 16918
rect 10888 16794 10916 18906
rect 10980 18834 11008 19246
rect 10968 18828 11020 18834
rect 10968 18770 11020 18776
rect 10980 18426 11008 18770
rect 10968 18420 11020 18426
rect 10968 18362 11020 18368
rect 10980 18170 11008 18362
rect 11152 18284 11204 18290
rect 11152 18226 11204 18232
rect 10980 18142 11100 18170
rect 10968 18080 11020 18086
rect 10968 18022 11020 18028
rect 10980 17678 11008 18022
rect 10968 17672 11020 17678
rect 10968 17614 11020 17620
rect 10968 17264 11020 17270
rect 10968 17206 11020 17212
rect 10692 16788 10744 16794
rect 10692 16730 10744 16736
rect 10876 16788 10928 16794
rect 10876 16730 10928 16736
rect 10704 16574 10732 16730
rect 10784 16584 10836 16590
rect 10704 16546 10784 16574
rect 10784 16526 10836 16532
rect 10876 16516 10928 16522
rect 10876 16458 10928 16464
rect 10692 16448 10744 16454
rect 10692 16390 10744 16396
rect 10704 15910 10732 16390
rect 10888 15910 10916 16458
rect 10692 15904 10744 15910
rect 10692 15846 10744 15852
rect 10876 15904 10928 15910
rect 10876 15846 10928 15852
rect 10704 15366 10732 15846
rect 10888 15570 10916 15846
rect 10876 15564 10928 15570
rect 10876 15506 10928 15512
rect 10980 15473 11008 17206
rect 11072 17134 11100 18142
rect 11164 17882 11192 18226
rect 11152 17876 11204 17882
rect 11152 17818 11204 17824
rect 11060 17128 11112 17134
rect 11060 17070 11112 17076
rect 11072 16794 11100 17070
rect 11060 16788 11112 16794
rect 11060 16730 11112 16736
rect 11152 16516 11204 16522
rect 11152 16458 11204 16464
rect 11164 15978 11192 16458
rect 11256 16114 11284 19246
rect 11336 19236 11388 19242
rect 11336 19178 11388 19184
rect 11244 16108 11296 16114
rect 11244 16050 11296 16056
rect 11152 15972 11204 15978
rect 11152 15914 11204 15920
rect 10966 15464 11022 15473
rect 10966 15399 11022 15408
rect 10692 15360 10744 15366
rect 10692 15302 10744 15308
rect 11164 15162 11192 15914
rect 11244 15904 11296 15910
rect 11244 15846 11296 15852
rect 11256 15502 11284 15846
rect 11244 15496 11296 15502
rect 11244 15438 11296 15444
rect 11152 15156 11204 15162
rect 11152 15098 11204 15104
rect 10600 15088 10652 15094
rect 10600 15030 10652 15036
rect 9312 15020 9364 15026
rect 9312 14962 9364 14968
rect 11348 14822 11376 19178
rect 11428 18624 11480 18630
rect 11428 18566 11480 18572
rect 11612 18624 11664 18630
rect 11612 18566 11664 18572
rect 11440 18426 11468 18566
rect 11428 18420 11480 18426
rect 11428 18362 11480 18368
rect 11520 18216 11572 18222
rect 11520 18158 11572 18164
rect 11532 17134 11560 18158
rect 11624 17270 11652 18566
rect 11980 17672 12032 17678
rect 11980 17614 12032 17620
rect 11612 17264 11664 17270
rect 11612 17206 11664 17212
rect 11520 17128 11572 17134
rect 11520 17070 11572 17076
rect 11888 16992 11940 16998
rect 11888 16934 11940 16940
rect 11900 16522 11928 16934
rect 11888 16516 11940 16522
rect 11888 16458 11940 16464
rect 11900 16250 11928 16458
rect 11992 16250 12020 17614
rect 12176 16794 12204 24822
rect 14740 24812 14792 24818
rect 14740 24754 14792 24760
rect 14648 24608 14700 24614
rect 14648 24550 14700 24556
rect 14660 24206 14688 24550
rect 12900 24200 12952 24206
rect 12900 24142 12952 24148
rect 14648 24200 14700 24206
rect 14648 24142 14700 24148
rect 12624 23112 12676 23118
rect 12624 23054 12676 23060
rect 12636 22778 12664 23054
rect 12624 22772 12676 22778
rect 12624 22714 12676 22720
rect 12532 22704 12584 22710
rect 12532 22646 12584 22652
rect 12440 22024 12492 22030
rect 12440 21966 12492 21972
rect 12348 21480 12400 21486
rect 12348 21422 12400 21428
rect 12360 20398 12388 21422
rect 12452 20942 12480 21966
rect 12544 21486 12572 22646
rect 12912 22642 12940 24142
rect 14752 23866 14780 24754
rect 14846 24508 15154 24528
rect 14846 24506 14852 24508
rect 14908 24506 14932 24508
rect 14988 24506 15012 24508
rect 15068 24506 15092 24508
rect 15148 24506 15154 24508
rect 14908 24454 14910 24506
rect 15090 24454 15092 24506
rect 14846 24452 14852 24454
rect 14908 24452 14932 24454
rect 14988 24452 15012 24454
rect 15068 24452 15092 24454
rect 15148 24452 15154 24454
rect 14846 24432 15154 24452
rect 16304 24200 16356 24206
rect 16304 24142 16356 24148
rect 15568 24064 15620 24070
rect 15568 24006 15620 24012
rect 14740 23860 14792 23866
rect 14740 23802 14792 23808
rect 15292 23792 15344 23798
rect 15292 23734 15344 23740
rect 14846 23420 15154 23440
rect 14846 23418 14852 23420
rect 14908 23418 14932 23420
rect 14988 23418 15012 23420
rect 15068 23418 15092 23420
rect 15148 23418 15154 23420
rect 14908 23366 14910 23418
rect 15090 23366 15092 23418
rect 14846 23364 14852 23366
rect 14908 23364 14932 23366
rect 14988 23364 15012 23366
rect 15068 23364 15092 23366
rect 15148 23364 15154 23366
rect 14846 23344 15154 23364
rect 15304 23322 15332 23734
rect 15580 23730 15608 24006
rect 16316 23866 16344 24142
rect 16396 24064 16448 24070
rect 16396 24006 16448 24012
rect 16948 24064 17000 24070
rect 16948 24006 17000 24012
rect 17224 24064 17276 24070
rect 17224 24006 17276 24012
rect 16408 23866 16436 24006
rect 16304 23860 16356 23866
rect 16304 23802 16356 23808
rect 16396 23860 16448 23866
rect 16396 23802 16448 23808
rect 16960 23730 16988 24006
rect 17132 23792 17184 23798
rect 17132 23734 17184 23740
rect 15568 23724 15620 23730
rect 15568 23666 15620 23672
rect 16120 23724 16172 23730
rect 16120 23666 16172 23672
rect 16948 23724 17000 23730
rect 16948 23666 17000 23672
rect 15476 23656 15528 23662
rect 15476 23598 15528 23604
rect 15292 23316 15344 23322
rect 15292 23258 15344 23264
rect 13452 23112 13504 23118
rect 13452 23054 13504 23060
rect 12992 22976 13044 22982
rect 12992 22918 13044 22924
rect 13268 22976 13320 22982
rect 13268 22918 13320 22924
rect 13004 22710 13032 22918
rect 12992 22704 13044 22710
rect 12992 22646 13044 22652
rect 12900 22636 12952 22642
rect 12900 22578 12952 22584
rect 12912 22030 12940 22578
rect 12900 22024 12952 22030
rect 12900 21966 12952 21972
rect 13280 21962 13308 22918
rect 13268 21956 13320 21962
rect 13268 21898 13320 21904
rect 12716 21888 12768 21894
rect 12636 21836 12716 21842
rect 12636 21830 12768 21836
rect 12636 21814 12756 21830
rect 12636 21622 12664 21814
rect 13464 21690 13492 23054
rect 15304 22710 15332 23258
rect 15488 23254 15516 23598
rect 15476 23248 15528 23254
rect 15476 23190 15528 23196
rect 15580 22982 15608 23666
rect 15660 23520 15712 23526
rect 15660 23462 15712 23468
rect 15672 23186 15700 23462
rect 16132 23322 16160 23666
rect 17040 23520 17092 23526
rect 17040 23462 17092 23468
rect 16120 23316 16172 23322
rect 16120 23258 16172 23264
rect 16488 23248 16540 23254
rect 16488 23190 16540 23196
rect 15660 23180 15712 23186
rect 15660 23122 15712 23128
rect 15568 22976 15620 22982
rect 15568 22918 15620 22924
rect 15292 22704 15344 22710
rect 15292 22646 15344 22652
rect 14188 22568 14240 22574
rect 14188 22510 14240 22516
rect 13912 22500 13964 22506
rect 13912 22442 13964 22448
rect 13924 21894 13952 22442
rect 13912 21888 13964 21894
rect 13912 21830 13964 21836
rect 14004 21888 14056 21894
rect 14004 21830 14056 21836
rect 13924 21690 13952 21830
rect 13452 21684 13504 21690
rect 13452 21626 13504 21632
rect 13912 21684 13964 21690
rect 13912 21626 13964 21632
rect 12624 21616 12676 21622
rect 12624 21558 12676 21564
rect 12532 21480 12584 21486
rect 12532 21422 12584 21428
rect 12440 20936 12492 20942
rect 12440 20878 12492 20884
rect 12348 20392 12400 20398
rect 12348 20334 12400 20340
rect 12360 20058 12388 20334
rect 12348 20052 12400 20058
rect 12348 19994 12400 20000
rect 12256 19712 12308 19718
rect 12256 19654 12308 19660
rect 12268 19446 12296 19654
rect 12256 19440 12308 19446
rect 12256 19382 12308 19388
rect 12268 18698 12296 19382
rect 12256 18692 12308 18698
rect 12256 18634 12308 18640
rect 12360 17270 12388 19994
rect 12544 19378 12572 21422
rect 12532 19372 12584 19378
rect 12532 19314 12584 19320
rect 12440 18624 12492 18630
rect 12440 18566 12492 18572
rect 12452 17542 12480 18566
rect 12636 17610 12664 21558
rect 14016 21554 14044 21830
rect 14004 21548 14056 21554
rect 14004 21490 14056 21496
rect 13452 21344 13504 21350
rect 13452 21286 13504 21292
rect 13464 20806 13492 21286
rect 13544 20936 13596 20942
rect 13544 20878 13596 20884
rect 12808 20800 12860 20806
rect 12808 20742 12860 20748
rect 13452 20800 13504 20806
rect 13452 20742 13504 20748
rect 12820 20466 12848 20742
rect 12808 20460 12860 20466
rect 12808 20402 12860 20408
rect 12716 18964 12768 18970
rect 12716 18906 12768 18912
rect 12728 17882 12756 18906
rect 12820 18698 12848 20402
rect 13084 19848 13136 19854
rect 13084 19790 13136 19796
rect 13096 19310 13124 19790
rect 13084 19304 13136 19310
rect 13084 19246 13136 19252
rect 12808 18692 12860 18698
rect 12808 18634 12860 18640
rect 13096 18358 13124 19246
rect 13084 18352 13136 18358
rect 13084 18294 13136 18300
rect 13360 18080 13412 18086
rect 13360 18022 13412 18028
rect 13372 17882 13400 18022
rect 12716 17876 12768 17882
rect 12716 17818 12768 17824
rect 13360 17876 13412 17882
rect 13360 17818 13412 17824
rect 12992 17808 13044 17814
rect 12992 17750 13044 17756
rect 12808 17672 12860 17678
rect 12808 17614 12860 17620
rect 12624 17604 12676 17610
rect 12624 17546 12676 17552
rect 12440 17536 12492 17542
rect 12440 17478 12492 17484
rect 12348 17264 12400 17270
rect 12348 17206 12400 17212
rect 12256 17196 12308 17202
rect 12256 17138 12308 17144
rect 12164 16788 12216 16794
rect 12164 16730 12216 16736
rect 11888 16244 11940 16250
rect 11888 16186 11940 16192
rect 11980 16244 12032 16250
rect 11980 16186 12032 16192
rect 11428 16108 11480 16114
rect 11428 16050 11480 16056
rect 11704 16108 11756 16114
rect 11704 16050 11756 16056
rect 11440 15026 11468 16050
rect 11716 15706 11744 16050
rect 11900 15706 11928 16186
rect 12268 16046 12296 17138
rect 12714 17096 12770 17105
rect 12714 17031 12770 17040
rect 12256 16040 12308 16046
rect 12256 15982 12308 15988
rect 11704 15700 11756 15706
rect 11704 15642 11756 15648
rect 11888 15700 11940 15706
rect 11888 15642 11940 15648
rect 12348 15428 12400 15434
rect 12348 15370 12400 15376
rect 12532 15428 12584 15434
rect 12532 15370 12584 15376
rect 12360 15026 12388 15370
rect 12544 15162 12572 15370
rect 12532 15156 12584 15162
rect 12532 15098 12584 15104
rect 11428 15020 11480 15026
rect 11428 14962 11480 14968
rect 11980 15020 12032 15026
rect 11980 14962 12032 14968
rect 12348 15020 12400 15026
rect 12348 14962 12400 14968
rect 9404 14816 9456 14822
rect 9404 14758 9456 14764
rect 11336 14816 11388 14822
rect 11336 14758 11388 14764
rect 8668 14544 8720 14550
rect 8668 14486 8720 14492
rect 8300 14408 8352 14414
rect 8300 14350 8352 14356
rect 8312 13870 8340 14350
rect 8484 14272 8536 14278
rect 8484 14214 8536 14220
rect 8496 13938 8524 14214
rect 8484 13932 8536 13938
rect 8484 13874 8536 13880
rect 8576 13932 8628 13938
rect 8576 13874 8628 13880
rect 8300 13864 8352 13870
rect 8300 13806 8352 13812
rect 8208 13728 8260 13734
rect 8208 13670 8260 13676
rect 8116 13524 8168 13530
rect 8116 13466 8168 13472
rect 8220 13462 8248 13670
rect 8208 13456 8260 13462
rect 8208 13398 8260 13404
rect 8208 13184 8260 13190
rect 8208 13126 8260 13132
rect 8024 12776 8076 12782
rect 8076 12724 8156 12730
rect 8024 12718 8156 12724
rect 8036 12702 8156 12718
rect 8128 12374 8156 12702
rect 8220 12646 8248 13126
rect 8208 12640 8260 12646
rect 8208 12582 8260 12588
rect 8024 12368 8076 12374
rect 8024 12310 8076 12316
rect 8116 12368 8168 12374
rect 8116 12310 8168 12316
rect 8036 12102 8064 12310
rect 7748 12096 7800 12102
rect 7748 12038 7800 12044
rect 8024 12096 8076 12102
rect 8024 12038 8076 12044
rect 7656 11756 7708 11762
rect 7656 11698 7708 11704
rect 7564 11688 7616 11694
rect 7392 11614 7512 11642
rect 7564 11630 7616 11636
rect 7484 10674 7512 11614
rect 7472 10668 7524 10674
rect 7472 10610 7524 10616
rect 7288 10260 7340 10266
rect 7288 10202 7340 10208
rect 7104 10056 7156 10062
rect 7104 9998 7156 10004
rect 6920 9444 6972 9450
rect 6920 9386 6972 9392
rect 7116 9382 7144 9998
rect 7484 9625 7512 10610
rect 7576 10470 7604 11630
rect 7656 11620 7708 11626
rect 7656 11562 7708 11568
rect 7668 11286 7696 11562
rect 7656 11280 7708 11286
rect 7656 11222 7708 11228
rect 7760 11150 7788 12038
rect 7840 11892 7892 11898
rect 7840 11834 7892 11840
rect 7748 11144 7800 11150
rect 7748 11086 7800 11092
rect 7852 10810 7880 11834
rect 8128 11150 8156 12310
rect 8208 12164 8260 12170
rect 8208 12106 8260 12112
rect 8220 11694 8248 12106
rect 8208 11688 8260 11694
rect 8208 11630 8260 11636
rect 8220 11150 8248 11630
rect 8116 11144 8168 11150
rect 8116 11086 8168 11092
rect 8208 11144 8260 11150
rect 8208 11086 8260 11092
rect 8312 11082 8340 13806
rect 8392 13728 8444 13734
rect 8392 13670 8444 13676
rect 8404 13394 8432 13670
rect 8392 13388 8444 13394
rect 8392 13330 8444 13336
rect 8484 13252 8536 13258
rect 8484 13194 8536 13200
rect 8496 12850 8524 13194
rect 8484 12844 8536 12850
rect 8404 12804 8484 12832
rect 8404 12442 8432 12804
rect 8484 12786 8536 12792
rect 8588 12442 8616 13874
rect 8680 12782 8708 14486
rect 9416 14414 9444 14758
rect 9404 14408 9456 14414
rect 9404 14350 9456 14356
rect 8944 13932 8996 13938
rect 8944 13874 8996 13880
rect 8760 13252 8812 13258
rect 8760 13194 8812 13200
rect 8772 12986 8800 13194
rect 8956 13190 8984 13874
rect 9128 13728 9180 13734
rect 9128 13670 9180 13676
rect 9140 13326 9168 13670
rect 9416 13444 9444 14350
rect 9496 14272 9548 14278
rect 9496 14214 9548 14220
rect 9508 13734 9536 14214
rect 10214 14172 10522 14192
rect 10214 14170 10220 14172
rect 10276 14170 10300 14172
rect 10356 14170 10380 14172
rect 10436 14170 10460 14172
rect 10516 14170 10522 14172
rect 10276 14118 10278 14170
rect 10458 14118 10460 14170
rect 10214 14116 10220 14118
rect 10276 14116 10300 14118
rect 10356 14116 10380 14118
rect 10436 14116 10460 14118
rect 10516 14116 10522 14118
rect 10214 14096 10522 14116
rect 10140 14000 10192 14006
rect 10140 13942 10192 13948
rect 9588 13932 9640 13938
rect 9588 13874 9640 13880
rect 9496 13728 9548 13734
rect 9494 13696 9496 13705
rect 9548 13696 9550 13705
rect 9494 13631 9550 13640
rect 9508 13605 9536 13631
rect 9600 13530 9628 13874
rect 9588 13524 9640 13530
rect 9588 13466 9640 13472
rect 9496 13456 9548 13462
rect 9416 13416 9496 13444
rect 9496 13398 9548 13404
rect 9128 13320 9180 13326
rect 9128 13262 9180 13268
rect 8852 13184 8904 13190
rect 8852 13126 8904 13132
rect 8944 13184 8996 13190
rect 8944 13126 8996 13132
rect 8760 12980 8812 12986
rect 8760 12922 8812 12928
rect 8668 12776 8720 12782
rect 8668 12718 8720 12724
rect 8392 12436 8444 12442
rect 8392 12378 8444 12384
rect 8576 12436 8628 12442
rect 8576 12378 8628 12384
rect 8404 11762 8432 12378
rect 8668 12096 8720 12102
rect 8668 12038 8720 12044
rect 8392 11756 8444 11762
rect 8392 11698 8444 11704
rect 8300 11076 8352 11082
rect 8300 11018 8352 11024
rect 7840 10804 7892 10810
rect 7840 10746 7892 10752
rect 8116 10804 8168 10810
rect 8116 10746 8168 10752
rect 7748 10668 7800 10674
rect 7748 10610 7800 10616
rect 7564 10464 7616 10470
rect 7564 10406 7616 10412
rect 7760 10130 7788 10610
rect 7748 10124 7800 10130
rect 7748 10066 7800 10072
rect 7760 9654 7788 10066
rect 7748 9648 7800 9654
rect 7470 9616 7526 9625
rect 7380 9580 7432 9586
rect 7748 9590 7800 9596
rect 7470 9551 7526 9560
rect 8024 9580 8076 9586
rect 7380 9522 7432 9528
rect 8024 9522 8076 9528
rect 6000 9376 6052 9382
rect 6000 9318 6052 9324
rect 7104 9376 7156 9382
rect 7104 9318 7156 9324
rect 5582 9276 5890 9296
rect 5582 9274 5588 9276
rect 5644 9274 5668 9276
rect 5724 9274 5748 9276
rect 5804 9274 5828 9276
rect 5884 9274 5890 9276
rect 5644 9222 5646 9274
rect 5826 9222 5828 9274
rect 5582 9220 5588 9222
rect 5644 9220 5668 9222
rect 5724 9220 5748 9222
rect 5804 9220 5828 9222
rect 5884 9220 5890 9222
rect 5582 9200 5890 9220
rect 1860 8968 1912 8974
rect 1858 8936 1860 8945
rect 4620 8968 4672 8974
rect 1912 8936 1914 8945
rect 4620 8910 4672 8916
rect 1858 8871 1914 8880
rect 4632 8430 4660 8910
rect 6828 8900 6880 8906
rect 6828 8842 6880 8848
rect 6840 8634 6868 8842
rect 6828 8628 6880 8634
rect 6828 8570 6880 8576
rect 7116 8498 7144 9318
rect 7392 9178 7420 9522
rect 8036 9382 8064 9522
rect 8024 9376 8076 9382
rect 8024 9318 8076 9324
rect 7380 9172 7432 9178
rect 7380 9114 7432 9120
rect 8036 9110 8064 9318
rect 8024 9104 8076 9110
rect 8024 9046 8076 9052
rect 7932 8968 7984 8974
rect 7932 8910 7984 8916
rect 7656 8832 7708 8838
rect 7656 8774 7708 8780
rect 6368 8492 6420 8498
rect 6368 8434 6420 8440
rect 7104 8492 7156 8498
rect 7104 8434 7156 8440
rect 4620 8424 4672 8430
rect 1766 8392 1822 8401
rect 4620 8366 4672 8372
rect 1766 8327 1822 8336
rect 1398 8256 1454 8265
rect 1398 8191 1454 8200
rect 1412 8090 1440 8191
rect 1400 8084 1452 8090
rect 1400 8026 1452 8032
rect 4632 7410 4660 8366
rect 6092 8288 6144 8294
rect 6092 8230 6144 8236
rect 5582 8188 5890 8208
rect 5582 8186 5588 8188
rect 5644 8186 5668 8188
rect 5724 8186 5748 8188
rect 5804 8186 5828 8188
rect 5884 8186 5890 8188
rect 5644 8134 5646 8186
rect 5826 8134 5828 8186
rect 5582 8132 5588 8134
rect 5644 8132 5668 8134
rect 5724 8132 5748 8134
rect 5804 8132 5828 8134
rect 5884 8132 5890 8134
rect 5582 8112 5890 8132
rect 6104 7954 6132 8230
rect 6380 8090 6408 8434
rect 7668 8430 7696 8774
rect 7944 8498 7972 8910
rect 7932 8492 7984 8498
rect 7932 8434 7984 8440
rect 7656 8424 7708 8430
rect 7656 8366 7708 8372
rect 6920 8288 6972 8294
rect 6920 8230 6972 8236
rect 7656 8288 7708 8294
rect 7656 8230 7708 8236
rect 6368 8084 6420 8090
rect 6368 8026 6420 8032
rect 6092 7948 6144 7954
rect 6092 7890 6144 7896
rect 6932 7886 6960 8230
rect 7012 8016 7064 8022
rect 7012 7958 7064 7964
rect 7024 7886 7052 7958
rect 5908 7880 5960 7886
rect 5908 7822 5960 7828
rect 6920 7880 6972 7886
rect 6920 7822 6972 7828
rect 7012 7880 7064 7886
rect 7012 7822 7064 7828
rect 7564 7880 7616 7886
rect 7564 7822 7616 7828
rect 4620 7404 4672 7410
rect 4620 7346 4672 7352
rect 4632 6934 4660 7346
rect 5582 7100 5890 7120
rect 5582 7098 5588 7100
rect 5644 7098 5668 7100
rect 5724 7098 5748 7100
rect 5804 7098 5828 7100
rect 5884 7098 5890 7100
rect 5644 7046 5646 7098
rect 5826 7046 5828 7098
rect 5582 7044 5588 7046
rect 5644 7044 5668 7046
rect 5724 7044 5748 7046
rect 5804 7044 5828 7046
rect 5884 7044 5890 7046
rect 5582 7024 5890 7044
rect 5920 7002 5948 7822
rect 6460 7812 6512 7818
rect 6460 7754 6512 7760
rect 6644 7812 6696 7818
rect 6644 7754 6696 7760
rect 6736 7812 6788 7818
rect 6736 7754 6788 7760
rect 6472 7342 6500 7754
rect 6460 7336 6512 7342
rect 6460 7278 6512 7284
rect 5908 6996 5960 7002
rect 5908 6938 5960 6944
rect 4620 6928 4672 6934
rect 4620 6870 4672 6876
rect 5920 6662 5948 6938
rect 6368 6724 6420 6730
rect 6368 6666 6420 6672
rect 5908 6656 5960 6662
rect 5908 6598 5960 6604
rect 6380 6458 6408 6666
rect 6656 6458 6684 7754
rect 6748 7698 6776 7754
rect 7024 7698 7052 7822
rect 6748 7670 6868 7698
rect 6368 6452 6420 6458
rect 6368 6394 6420 6400
rect 6644 6452 6696 6458
rect 6644 6394 6696 6400
rect 6840 6322 6868 7670
rect 6932 7670 7052 7698
rect 6932 6798 6960 7670
rect 7012 7404 7064 7410
rect 7012 7346 7064 7352
rect 7024 6798 7052 7346
rect 7576 7342 7604 7822
rect 7668 7410 7696 8230
rect 7840 7880 7892 7886
rect 7944 7834 7972 8434
rect 8036 7886 8064 9046
rect 8128 8974 8156 10746
rect 8404 10266 8432 11698
rect 8680 10674 8708 12038
rect 8772 11694 8800 12922
rect 8864 12306 8892 13126
rect 8956 12918 8984 13126
rect 9508 12986 9536 13398
rect 9496 12980 9548 12986
rect 9496 12922 9548 12928
rect 8944 12912 8996 12918
rect 8944 12854 8996 12860
rect 9680 12776 9732 12782
rect 9680 12718 9732 12724
rect 9864 12776 9916 12782
rect 9864 12718 9916 12724
rect 9692 12442 9720 12718
rect 9680 12436 9732 12442
rect 9680 12378 9732 12384
rect 9876 12374 9904 12718
rect 9864 12368 9916 12374
rect 9864 12310 9916 12316
rect 10048 12368 10100 12374
rect 10048 12310 10100 12316
rect 8852 12300 8904 12306
rect 8852 12242 8904 12248
rect 8760 11688 8812 11694
rect 8760 11630 8812 11636
rect 8864 11150 8892 12242
rect 9680 12232 9732 12238
rect 9680 12174 9732 12180
rect 9312 12164 9364 12170
rect 9312 12106 9364 12112
rect 9324 11354 9352 12106
rect 9692 11762 9720 12174
rect 9680 11756 9732 11762
rect 9680 11698 9732 11704
rect 9312 11348 9364 11354
rect 9312 11290 9364 11296
rect 8852 11144 8904 11150
rect 8852 11086 8904 11092
rect 9496 11144 9548 11150
rect 9496 11086 9548 11092
rect 8944 11076 8996 11082
rect 8944 11018 8996 11024
rect 8956 10674 8984 11018
rect 8668 10668 8720 10674
rect 8668 10610 8720 10616
rect 8944 10668 8996 10674
rect 8944 10610 8996 10616
rect 8392 10260 8444 10266
rect 8392 10202 8444 10208
rect 8300 10056 8352 10062
rect 8300 9998 8352 10004
rect 8312 9654 8340 9998
rect 8300 9648 8352 9654
rect 8300 9590 8352 9596
rect 8116 8968 8168 8974
rect 8116 8910 8168 8916
rect 7892 7828 7972 7834
rect 7840 7822 7972 7828
rect 8024 7880 8076 7886
rect 8024 7822 8076 7828
rect 7852 7806 7972 7822
rect 7840 7744 7892 7750
rect 7840 7686 7892 7692
rect 7852 7478 7880 7686
rect 7840 7472 7892 7478
rect 7840 7414 7892 7420
rect 7656 7404 7708 7410
rect 7656 7346 7708 7352
rect 7564 7336 7616 7342
rect 7564 7278 7616 7284
rect 7104 6996 7156 7002
rect 7104 6938 7156 6944
rect 6920 6792 6972 6798
rect 6920 6734 6972 6740
rect 7012 6792 7064 6798
rect 7012 6734 7064 6740
rect 7116 6322 7144 6938
rect 7576 6322 7604 7278
rect 7944 6934 7972 7806
rect 8036 7002 8064 7822
rect 8116 7540 8168 7546
rect 8116 7482 8168 7488
rect 8024 6996 8076 7002
rect 8024 6938 8076 6944
rect 7932 6928 7984 6934
rect 7932 6870 7984 6876
rect 7944 6798 7972 6870
rect 7932 6792 7984 6798
rect 7932 6734 7984 6740
rect 7748 6656 7800 6662
rect 7748 6598 7800 6604
rect 7760 6390 7788 6598
rect 8128 6458 8156 7482
rect 8312 6662 8340 9590
rect 8680 9586 8892 9602
rect 8668 9580 8892 9586
rect 8720 9574 8892 9580
rect 8668 9522 8720 9528
rect 8864 9518 8892 9574
rect 8956 9518 8984 10610
rect 9036 10464 9088 10470
rect 9036 10406 9088 10412
rect 9048 10266 9076 10406
rect 9036 10260 9088 10266
rect 9036 10202 9088 10208
rect 9128 10124 9180 10130
rect 9128 10066 9180 10072
rect 9140 9722 9168 10066
rect 9220 10056 9272 10062
rect 9220 9998 9272 10004
rect 9312 10056 9364 10062
rect 9312 9998 9364 10004
rect 9128 9716 9180 9722
rect 9128 9658 9180 9664
rect 9126 9616 9182 9625
rect 9036 9580 9088 9586
rect 9126 9551 9128 9560
rect 9036 9522 9088 9528
rect 9180 9551 9182 9560
rect 9128 9522 9180 9528
rect 8852 9512 8904 9518
rect 8852 9454 8904 9460
rect 8944 9512 8996 9518
rect 8944 9454 8996 9460
rect 8484 9376 8536 9382
rect 8484 9318 8536 9324
rect 8668 9376 8720 9382
rect 9048 9364 9076 9522
rect 8720 9336 9076 9364
rect 8668 9318 8720 9324
rect 8496 9178 8524 9318
rect 9232 9178 9260 9998
rect 9324 9654 9352 9998
rect 9312 9648 9364 9654
rect 9312 9590 9364 9596
rect 8484 9172 8536 9178
rect 8484 9114 8536 9120
rect 9220 9172 9272 9178
rect 9220 9114 9272 9120
rect 8392 8900 8444 8906
rect 8392 8842 8444 8848
rect 8576 8900 8628 8906
rect 8576 8842 8628 8848
rect 8404 8498 8432 8842
rect 8484 8628 8536 8634
rect 8484 8570 8536 8576
rect 8392 8492 8444 8498
rect 8392 8434 8444 8440
rect 8404 7002 8432 8434
rect 8496 7410 8524 8570
rect 8588 8566 8616 8842
rect 8576 8560 8628 8566
rect 8576 8502 8628 8508
rect 8484 7404 8536 7410
rect 8484 7346 8536 7352
rect 8392 6996 8444 7002
rect 8392 6938 8444 6944
rect 8392 6792 8444 6798
rect 8392 6734 8444 6740
rect 8300 6656 8352 6662
rect 8300 6598 8352 6604
rect 8116 6452 8168 6458
rect 8116 6394 8168 6400
rect 7748 6384 7800 6390
rect 7748 6326 7800 6332
rect 6828 6316 6880 6322
rect 6828 6258 6880 6264
rect 7104 6316 7156 6322
rect 7104 6258 7156 6264
rect 7564 6316 7616 6322
rect 7564 6258 7616 6264
rect 7576 6118 7604 6258
rect 8312 6254 8340 6598
rect 8404 6458 8432 6734
rect 8496 6458 8524 7346
rect 9128 7268 9180 7274
rect 9128 7210 9180 7216
rect 9140 7002 9168 7210
rect 9232 7002 9260 9114
rect 9508 8634 9536 11086
rect 9692 10742 9720 11698
rect 9772 11552 9824 11558
rect 9772 11494 9824 11500
rect 9784 11354 9812 11494
rect 9772 11348 9824 11354
rect 9772 11290 9824 11296
rect 9876 11150 9904 12310
rect 10060 11762 10088 12310
rect 10048 11756 10100 11762
rect 10048 11698 10100 11704
rect 10152 11558 10180 13942
rect 10232 13728 10284 13734
rect 10232 13670 10284 13676
rect 10244 13258 10272 13670
rect 10232 13252 10284 13258
rect 10232 13194 10284 13200
rect 11152 13184 11204 13190
rect 11152 13126 11204 13132
rect 10214 13084 10522 13104
rect 10214 13082 10220 13084
rect 10276 13082 10300 13084
rect 10356 13082 10380 13084
rect 10436 13082 10460 13084
rect 10516 13082 10522 13084
rect 10276 13030 10278 13082
rect 10458 13030 10460 13082
rect 10214 13028 10220 13030
rect 10276 13028 10300 13030
rect 10356 13028 10380 13030
rect 10436 13028 10460 13030
rect 10516 13028 10522 13030
rect 10214 13008 10522 13028
rect 10968 12640 11020 12646
rect 10968 12582 11020 12588
rect 10600 12436 10652 12442
rect 10600 12378 10652 12384
rect 10214 11996 10522 12016
rect 10214 11994 10220 11996
rect 10276 11994 10300 11996
rect 10356 11994 10380 11996
rect 10436 11994 10460 11996
rect 10516 11994 10522 11996
rect 10276 11942 10278 11994
rect 10458 11942 10460 11994
rect 10214 11940 10220 11942
rect 10276 11940 10300 11942
rect 10356 11940 10380 11942
rect 10436 11940 10460 11942
rect 10516 11940 10522 11942
rect 10214 11920 10522 11940
rect 10230 11792 10286 11801
rect 10612 11762 10640 12378
rect 10876 12164 10928 12170
rect 10876 12106 10928 12112
rect 10888 11898 10916 12106
rect 10692 11892 10744 11898
rect 10692 11834 10744 11840
rect 10876 11892 10928 11898
rect 10876 11834 10928 11840
rect 10230 11727 10232 11736
rect 10284 11727 10286 11736
rect 10324 11756 10376 11762
rect 10232 11698 10284 11704
rect 10600 11756 10652 11762
rect 10376 11716 10456 11744
rect 10324 11698 10376 11704
rect 10324 11620 10376 11626
rect 10324 11562 10376 11568
rect 10140 11552 10192 11558
rect 10140 11494 10192 11500
rect 9864 11144 9916 11150
rect 9864 11086 9916 11092
rect 10152 11082 10180 11494
rect 10336 11257 10364 11562
rect 10428 11354 10456 11716
rect 10600 11698 10652 11704
rect 10600 11552 10652 11558
rect 10600 11494 10652 11500
rect 10416 11348 10468 11354
rect 10416 11290 10468 11296
rect 10322 11248 10378 11257
rect 10322 11183 10378 11192
rect 10612 11150 10640 11494
rect 10704 11286 10732 11834
rect 10980 11801 11008 12582
rect 11164 12238 11192 13126
rect 11152 12232 11204 12238
rect 11152 12174 11204 12180
rect 11164 11898 11192 12174
rect 11152 11892 11204 11898
rect 11152 11834 11204 11840
rect 10966 11792 11022 11801
rect 10966 11727 11022 11736
rect 10692 11280 10744 11286
rect 10692 11222 10744 11228
rect 10600 11144 10652 11150
rect 10600 11086 10652 11092
rect 10784 11144 10836 11150
rect 10968 11144 11020 11150
rect 10836 11092 10916 11098
rect 10784 11086 10916 11092
rect 10968 11086 11020 11092
rect 11150 11112 11206 11121
rect 10140 11076 10192 11082
rect 10796 11070 10916 11086
rect 10140 11018 10192 11024
rect 9680 10736 9732 10742
rect 9680 10678 9732 10684
rect 10152 10674 10180 11018
rect 10784 11008 10836 11014
rect 10784 10950 10836 10956
rect 10214 10908 10522 10928
rect 10214 10906 10220 10908
rect 10276 10906 10300 10908
rect 10356 10906 10380 10908
rect 10436 10906 10460 10908
rect 10516 10906 10522 10908
rect 10276 10854 10278 10906
rect 10458 10854 10460 10906
rect 10214 10852 10220 10854
rect 10276 10852 10300 10854
rect 10356 10852 10380 10854
rect 10436 10852 10460 10854
rect 10516 10852 10522 10854
rect 10214 10832 10522 10852
rect 10140 10668 10192 10674
rect 10140 10610 10192 10616
rect 10796 10198 10824 10950
rect 10888 10810 10916 11070
rect 10980 10810 11008 11086
rect 11150 11047 11152 11056
rect 11204 11047 11206 11056
rect 11152 11018 11204 11024
rect 11244 11008 11296 11014
rect 11244 10950 11296 10956
rect 10876 10804 10928 10810
rect 10876 10746 10928 10752
rect 10968 10804 11020 10810
rect 10968 10746 11020 10752
rect 11256 10742 11284 10950
rect 11244 10736 11296 10742
rect 11244 10678 11296 10684
rect 11152 10464 11204 10470
rect 11152 10406 11204 10412
rect 10784 10192 10836 10198
rect 10784 10134 10836 10140
rect 11164 10130 11192 10406
rect 11152 10124 11204 10130
rect 11152 10066 11204 10072
rect 10214 9820 10522 9840
rect 10214 9818 10220 9820
rect 10276 9818 10300 9820
rect 10356 9818 10380 9820
rect 10436 9818 10460 9820
rect 10516 9818 10522 9820
rect 10276 9766 10278 9818
rect 10458 9766 10460 9818
rect 10214 9764 10220 9766
rect 10276 9764 10300 9766
rect 10356 9764 10380 9766
rect 10436 9764 10460 9766
rect 10516 9764 10522 9766
rect 10214 9744 10522 9764
rect 11164 9654 11192 10066
rect 11152 9648 11204 9654
rect 11152 9590 11204 9596
rect 9772 9580 9824 9586
rect 9772 9522 9824 9528
rect 9784 9178 9812 9522
rect 10508 9512 10560 9518
rect 10508 9454 10560 9460
rect 9772 9172 9824 9178
rect 9772 9114 9824 9120
rect 10520 9042 10548 9454
rect 11152 9444 11204 9450
rect 11152 9386 11204 9392
rect 10876 9376 10928 9382
rect 10876 9318 10928 9324
rect 10048 9036 10100 9042
rect 10048 8978 10100 8984
rect 10508 9036 10560 9042
rect 10508 8978 10560 8984
rect 9496 8628 9548 8634
rect 9496 8570 9548 8576
rect 9678 8528 9734 8537
rect 9678 8463 9680 8472
rect 9732 8463 9734 8472
rect 9680 8434 9732 8440
rect 10060 8072 10088 8978
rect 10140 8832 10192 8838
rect 10140 8774 10192 8780
rect 10152 8634 10180 8774
rect 10214 8732 10522 8752
rect 10214 8730 10220 8732
rect 10276 8730 10300 8732
rect 10356 8730 10380 8732
rect 10436 8730 10460 8732
rect 10516 8730 10522 8732
rect 10276 8678 10278 8730
rect 10458 8678 10460 8730
rect 10214 8676 10220 8678
rect 10276 8676 10300 8678
rect 10356 8676 10380 8678
rect 10436 8676 10460 8678
rect 10516 8676 10522 8678
rect 10214 8656 10522 8676
rect 10140 8628 10192 8634
rect 10140 8570 10192 8576
rect 10692 8560 10744 8566
rect 10692 8502 10744 8508
rect 10416 8492 10468 8498
rect 10416 8434 10468 8440
rect 10600 8492 10652 8498
rect 10600 8434 10652 8440
rect 10428 8090 10456 8434
rect 10508 8356 10560 8362
rect 10508 8298 10560 8304
rect 10416 8084 10468 8090
rect 10060 8044 10180 8072
rect 10046 7984 10102 7993
rect 10046 7919 10102 7928
rect 10060 7886 10088 7919
rect 10048 7880 10100 7886
rect 10048 7822 10100 7828
rect 9864 7404 9916 7410
rect 9916 7364 9996 7392
rect 9864 7346 9916 7352
rect 9772 7268 9824 7274
rect 9772 7210 9824 7216
rect 8576 6996 8628 7002
rect 8576 6938 8628 6944
rect 9128 6996 9180 7002
rect 9128 6938 9180 6944
rect 9220 6996 9272 7002
rect 9220 6938 9272 6944
rect 8392 6452 8444 6458
rect 8392 6394 8444 6400
rect 8484 6452 8536 6458
rect 8484 6394 8536 6400
rect 8300 6248 8352 6254
rect 8300 6190 8352 6196
rect 8496 6186 8524 6394
rect 8484 6180 8536 6186
rect 8484 6122 8536 6128
rect 7564 6112 7616 6118
rect 7564 6054 7616 6060
rect 5582 6012 5890 6032
rect 5582 6010 5588 6012
rect 5644 6010 5668 6012
rect 5724 6010 5748 6012
rect 5804 6010 5828 6012
rect 5884 6010 5890 6012
rect 5644 5958 5646 6010
rect 5826 5958 5828 6010
rect 5582 5956 5588 5958
rect 5644 5956 5668 5958
rect 5724 5956 5748 5958
rect 5804 5956 5828 5958
rect 5884 5956 5890 5958
rect 5582 5936 5890 5956
rect 8482 5944 8538 5953
rect 8482 5879 8484 5888
rect 8536 5879 8538 5888
rect 8484 5850 8536 5856
rect 8116 5772 8168 5778
rect 8116 5714 8168 5720
rect 1492 5568 1544 5574
rect 1490 5536 1492 5545
rect 1544 5536 1546 5545
rect 1490 5471 1546 5480
rect 8128 5302 8156 5714
rect 8496 5710 8524 5850
rect 8588 5778 8616 6938
rect 9680 6724 9732 6730
rect 9680 6666 9732 6672
rect 9692 6186 9720 6666
rect 9784 6390 9812 7210
rect 9968 7206 9996 7364
rect 9864 7200 9916 7206
rect 9864 7142 9916 7148
rect 9956 7200 10008 7206
rect 9956 7142 10008 7148
rect 9876 6458 9904 7142
rect 9968 6458 9996 7142
rect 10048 6656 10100 6662
rect 10048 6598 10100 6604
rect 9864 6452 9916 6458
rect 9864 6394 9916 6400
rect 9956 6452 10008 6458
rect 9956 6394 10008 6400
rect 9772 6384 9824 6390
rect 9772 6326 9824 6332
rect 9864 6248 9916 6254
rect 9864 6190 9916 6196
rect 9680 6180 9732 6186
rect 9680 6122 9732 6128
rect 9680 5840 9732 5846
rect 9680 5782 9732 5788
rect 8576 5772 8628 5778
rect 8576 5714 8628 5720
rect 9312 5772 9364 5778
rect 9312 5714 9364 5720
rect 8484 5704 8536 5710
rect 8484 5646 8536 5652
rect 9324 5370 9352 5714
rect 9588 5568 9640 5574
rect 9588 5510 9640 5516
rect 9312 5364 9364 5370
rect 9312 5306 9364 5312
rect 8116 5296 8168 5302
rect 8116 5238 8168 5244
rect 5582 4924 5890 4944
rect 5582 4922 5588 4924
rect 5644 4922 5668 4924
rect 5724 4922 5748 4924
rect 5804 4922 5828 4924
rect 5884 4922 5890 4924
rect 5644 4870 5646 4922
rect 5826 4870 5828 4922
rect 5582 4868 5588 4870
rect 5644 4868 5668 4870
rect 5724 4868 5748 4870
rect 5804 4868 5828 4870
rect 5884 4868 5890 4870
rect 5582 4848 5890 4868
rect 8128 4146 8156 5238
rect 9324 4622 9352 5306
rect 9600 5234 9628 5510
rect 9692 5370 9720 5782
rect 9680 5364 9732 5370
rect 9680 5306 9732 5312
rect 9876 5302 9904 6190
rect 9968 5574 9996 6394
rect 10060 5710 10088 6598
rect 10152 6254 10180 8044
rect 10416 8026 10468 8032
rect 10520 7954 10548 8298
rect 10508 7948 10560 7954
rect 10508 7890 10560 7896
rect 10612 7886 10640 8434
rect 10704 8430 10732 8502
rect 10888 8498 10916 9318
rect 10968 9104 11020 9110
rect 10968 9046 11020 9052
rect 10876 8492 10928 8498
rect 10876 8434 10928 8440
rect 10692 8424 10744 8430
rect 10692 8366 10744 8372
rect 10704 8294 10732 8366
rect 10692 8288 10744 8294
rect 10692 8230 10744 8236
rect 10888 8090 10916 8434
rect 10876 8084 10928 8090
rect 10876 8026 10928 8032
rect 10600 7880 10652 7886
rect 10600 7822 10652 7828
rect 10214 7644 10522 7664
rect 10214 7642 10220 7644
rect 10276 7642 10300 7644
rect 10356 7642 10380 7644
rect 10436 7642 10460 7644
rect 10516 7642 10522 7644
rect 10276 7590 10278 7642
rect 10458 7590 10460 7642
rect 10214 7588 10220 7590
rect 10276 7588 10300 7590
rect 10356 7588 10380 7590
rect 10436 7588 10460 7590
rect 10516 7588 10522 7590
rect 10214 7568 10522 7588
rect 10508 7404 10560 7410
rect 10612 7392 10640 7822
rect 10692 7744 10744 7750
rect 10692 7686 10744 7692
rect 10560 7364 10640 7392
rect 10508 7346 10560 7352
rect 10520 7002 10548 7346
rect 10508 6996 10560 7002
rect 10508 6938 10560 6944
rect 10600 6656 10652 6662
rect 10600 6598 10652 6604
rect 10214 6556 10522 6576
rect 10214 6554 10220 6556
rect 10276 6554 10300 6556
rect 10356 6554 10380 6556
rect 10436 6554 10460 6556
rect 10516 6554 10522 6556
rect 10276 6502 10278 6554
rect 10458 6502 10460 6554
rect 10214 6500 10220 6502
rect 10276 6500 10300 6502
rect 10356 6500 10380 6502
rect 10436 6500 10460 6502
rect 10516 6500 10522 6502
rect 10214 6480 10522 6500
rect 10612 6322 10640 6598
rect 10600 6316 10652 6322
rect 10600 6258 10652 6264
rect 10140 6248 10192 6254
rect 10140 6190 10192 6196
rect 10704 5914 10732 7686
rect 10980 7546 11008 9046
rect 11060 7812 11112 7818
rect 11060 7754 11112 7760
rect 10968 7540 11020 7546
rect 10888 7500 10968 7528
rect 10784 7336 10836 7342
rect 10784 7278 10836 7284
rect 10796 6798 10824 7278
rect 10784 6792 10836 6798
rect 10784 6734 10836 6740
rect 10692 5908 10744 5914
rect 10692 5850 10744 5856
rect 10048 5704 10100 5710
rect 10048 5646 10100 5652
rect 10140 5704 10192 5710
rect 10600 5704 10652 5710
rect 10140 5646 10192 5652
rect 10598 5672 10600 5681
rect 10652 5672 10654 5681
rect 9956 5568 10008 5574
rect 9956 5510 10008 5516
rect 9864 5296 9916 5302
rect 9864 5238 9916 5244
rect 9588 5228 9640 5234
rect 9588 5170 9640 5176
rect 9956 5092 10008 5098
rect 9956 5034 10008 5040
rect 9312 4616 9364 4622
rect 9312 4558 9364 4564
rect 9968 4146 9996 5034
rect 10060 5030 10088 5646
rect 10152 5234 10180 5646
rect 10704 5658 10732 5850
rect 10784 5772 10836 5778
rect 10888 5760 10916 7500
rect 10968 7482 11020 7488
rect 11072 7478 11100 7754
rect 11164 7562 11192 9386
rect 11244 9376 11296 9382
rect 11244 9318 11296 9324
rect 11256 8294 11284 9318
rect 11244 8288 11296 8294
rect 11244 8230 11296 8236
rect 11164 7534 11284 7562
rect 11060 7472 11112 7478
rect 11060 7414 11112 7420
rect 11072 6390 11100 7414
rect 11152 7404 11204 7410
rect 11152 7346 11204 7352
rect 11164 6798 11192 7346
rect 11152 6792 11204 6798
rect 11152 6734 11204 6740
rect 11060 6384 11112 6390
rect 11060 6326 11112 6332
rect 10836 5732 10916 5760
rect 10784 5714 10836 5720
rect 10704 5630 10824 5658
rect 10598 5607 10654 5616
rect 10692 5568 10744 5574
rect 10692 5510 10744 5516
rect 10214 5468 10522 5488
rect 10214 5466 10220 5468
rect 10276 5466 10300 5468
rect 10356 5466 10380 5468
rect 10436 5466 10460 5468
rect 10516 5466 10522 5468
rect 10276 5414 10278 5466
rect 10458 5414 10460 5466
rect 10214 5412 10220 5414
rect 10276 5412 10300 5414
rect 10356 5412 10380 5414
rect 10436 5412 10460 5414
rect 10516 5412 10522 5414
rect 10214 5392 10522 5412
rect 10704 5234 10732 5510
rect 10140 5228 10192 5234
rect 10140 5170 10192 5176
rect 10692 5228 10744 5234
rect 10692 5170 10744 5176
rect 10048 5024 10100 5030
rect 10048 4966 10100 4972
rect 10152 4826 10180 5170
rect 10416 5160 10468 5166
rect 10416 5102 10468 5108
rect 10140 4820 10192 4826
rect 10140 4762 10192 4768
rect 10140 4684 10192 4690
rect 10140 4626 10192 4632
rect 8116 4140 8168 4146
rect 8116 4082 8168 4088
rect 9956 4140 10008 4146
rect 9956 4082 10008 4088
rect 5582 3836 5890 3856
rect 5582 3834 5588 3836
rect 5644 3834 5668 3836
rect 5724 3834 5748 3836
rect 5804 3834 5828 3836
rect 5884 3834 5890 3836
rect 5644 3782 5646 3834
rect 5826 3782 5828 3834
rect 5582 3780 5588 3782
rect 5644 3780 5668 3782
rect 5724 3780 5748 3782
rect 5804 3780 5828 3782
rect 5884 3780 5890 3782
rect 5582 3760 5890 3780
rect 8128 3058 8156 4082
rect 10152 3942 10180 4626
rect 10428 4622 10456 5102
rect 10796 4622 10824 5630
rect 11060 5636 11112 5642
rect 11060 5578 11112 5584
rect 10876 5228 10928 5234
rect 10876 5170 10928 5176
rect 10416 4616 10468 4622
rect 10784 4616 10836 4622
rect 10468 4576 10640 4604
rect 10416 4558 10468 4564
rect 10214 4380 10522 4400
rect 10214 4378 10220 4380
rect 10276 4378 10300 4380
rect 10356 4378 10380 4380
rect 10436 4378 10460 4380
rect 10516 4378 10522 4380
rect 10276 4326 10278 4378
rect 10458 4326 10460 4378
rect 10214 4324 10220 4326
rect 10276 4324 10300 4326
rect 10356 4324 10380 4326
rect 10436 4324 10460 4326
rect 10516 4324 10522 4326
rect 10214 4304 10522 4324
rect 10612 4146 10640 4576
rect 10784 4558 10836 4564
rect 10600 4140 10652 4146
rect 10600 4082 10652 4088
rect 10796 4078 10824 4558
rect 10784 4072 10836 4078
rect 10784 4014 10836 4020
rect 10140 3936 10192 3942
rect 10140 3878 10192 3884
rect 10888 3534 10916 5170
rect 11072 5030 11100 5578
rect 11256 5370 11284 7534
rect 11348 6798 11376 14758
rect 11992 14618 12020 14962
rect 11980 14612 12032 14618
rect 11980 14554 12032 14560
rect 12624 14544 12676 14550
rect 12624 14486 12676 14492
rect 11980 14408 12032 14414
rect 11980 14350 12032 14356
rect 11704 13932 11756 13938
rect 11704 13874 11756 13880
rect 11716 13734 11744 13874
rect 11704 13728 11756 13734
rect 11704 13670 11756 13676
rect 11716 13394 11744 13670
rect 11704 13388 11756 13394
rect 11704 13330 11756 13336
rect 11612 12776 11664 12782
rect 11612 12718 11664 12724
rect 11624 12442 11652 12718
rect 11612 12436 11664 12442
rect 11612 12378 11664 12384
rect 11992 12306 12020 14350
rect 12440 14000 12492 14006
rect 12440 13942 12492 13948
rect 12164 13932 12216 13938
rect 12164 13874 12216 13880
rect 12176 13530 12204 13874
rect 12452 13802 12480 13942
rect 12532 13932 12584 13938
rect 12532 13874 12584 13880
rect 12440 13796 12492 13802
rect 12440 13738 12492 13744
rect 12164 13524 12216 13530
rect 12164 13466 12216 13472
rect 12072 13320 12124 13326
rect 12072 13262 12124 13268
rect 12084 12782 12112 13262
rect 12544 12986 12572 13874
rect 12636 13326 12664 14486
rect 12624 13320 12676 13326
rect 12624 13262 12676 13268
rect 12532 12980 12584 12986
rect 12532 12922 12584 12928
rect 12348 12912 12400 12918
rect 12348 12854 12400 12860
rect 12072 12776 12124 12782
rect 12072 12718 12124 12724
rect 12360 12442 12388 12854
rect 12728 12646 12756 17031
rect 12820 15910 12848 17614
rect 13004 17066 13032 17750
rect 13268 17332 13320 17338
rect 13268 17274 13320 17280
rect 12992 17060 13044 17066
rect 12992 17002 13044 17008
rect 13280 16998 13308 17274
rect 13268 16992 13320 16998
rect 13268 16934 13320 16940
rect 12900 16448 12952 16454
rect 12898 16416 12900 16425
rect 12952 16416 12954 16425
rect 12898 16351 12954 16360
rect 13280 16182 13308 16934
rect 13360 16584 13412 16590
rect 13358 16552 13360 16561
rect 13412 16552 13414 16561
rect 13358 16487 13414 16496
rect 13268 16176 13320 16182
rect 13268 16118 13320 16124
rect 13464 16028 13492 20742
rect 13556 20330 13584 20878
rect 13636 20460 13688 20466
rect 13636 20402 13688 20408
rect 13544 20324 13596 20330
rect 13544 20266 13596 20272
rect 13556 19922 13584 20266
rect 13544 19916 13596 19922
rect 13544 19858 13596 19864
rect 13648 19514 13676 20402
rect 13912 20256 13964 20262
rect 13912 20198 13964 20204
rect 13924 19854 13952 20198
rect 13912 19848 13964 19854
rect 13912 19790 13964 19796
rect 14016 19700 14044 21490
rect 14200 21486 14228 22510
rect 14846 22332 15154 22352
rect 14846 22330 14852 22332
rect 14908 22330 14932 22332
rect 14988 22330 15012 22332
rect 15068 22330 15092 22332
rect 15148 22330 15154 22332
rect 14908 22278 14910 22330
rect 15090 22278 15092 22330
rect 14846 22276 14852 22278
rect 14908 22276 14932 22278
rect 14988 22276 15012 22278
rect 15068 22276 15092 22278
rect 15148 22276 15154 22278
rect 14846 22256 15154 22276
rect 15580 22094 15608 22918
rect 15396 22066 15608 22094
rect 15672 22094 15700 23122
rect 15752 23112 15804 23118
rect 15752 23054 15804 23060
rect 15764 22234 15792 23054
rect 15844 22976 15896 22982
rect 15844 22918 15896 22924
rect 15856 22778 15884 22918
rect 15844 22772 15896 22778
rect 15844 22714 15896 22720
rect 15844 22636 15896 22642
rect 15844 22578 15896 22584
rect 15936 22636 15988 22642
rect 15936 22578 15988 22584
rect 15856 22506 15884 22578
rect 15844 22500 15896 22506
rect 15844 22442 15896 22448
rect 15752 22228 15804 22234
rect 15752 22170 15804 22176
rect 15948 22094 15976 22578
rect 16500 22166 16528 23190
rect 17052 22982 17080 23462
rect 17144 22982 17172 23734
rect 17236 23322 17264 24006
rect 17224 23316 17276 23322
rect 17224 23258 17276 23264
rect 17236 23118 17264 23258
rect 17224 23112 17276 23118
rect 17224 23054 17276 23060
rect 17040 22976 17092 22982
rect 17040 22918 17092 22924
rect 17132 22976 17184 22982
rect 17132 22918 17184 22924
rect 17960 22976 18012 22982
rect 17960 22918 18012 22924
rect 18236 22976 18288 22982
rect 18236 22918 18288 22924
rect 16672 22432 16724 22438
rect 16672 22374 16724 22380
rect 16684 22234 16712 22374
rect 16672 22228 16724 22234
rect 16672 22170 16724 22176
rect 16488 22160 16540 22166
rect 16488 22102 16540 22108
rect 15672 22066 15792 22094
rect 15292 21616 15344 21622
rect 15292 21558 15344 21564
rect 14188 21480 14240 21486
rect 14188 21422 14240 21428
rect 14846 21244 15154 21264
rect 14846 21242 14852 21244
rect 14908 21242 14932 21244
rect 14988 21242 15012 21244
rect 15068 21242 15092 21244
rect 15148 21242 15154 21244
rect 14908 21190 14910 21242
rect 15090 21190 15092 21242
rect 14846 21188 14852 21190
rect 14908 21188 14932 21190
rect 14988 21188 15012 21190
rect 15068 21188 15092 21190
rect 15148 21188 15154 21190
rect 14846 21168 15154 21188
rect 15304 20942 15332 21558
rect 15292 20936 15344 20942
rect 15292 20878 15344 20884
rect 14280 20460 14332 20466
rect 14280 20402 14332 20408
rect 14292 19718 14320 20402
rect 14556 20256 14608 20262
rect 14556 20198 14608 20204
rect 13924 19672 14044 19700
rect 14280 19712 14332 19718
rect 13636 19508 13688 19514
rect 13636 19450 13688 19456
rect 13820 18896 13872 18902
rect 13820 18838 13872 18844
rect 13832 18426 13860 18838
rect 13820 18420 13872 18426
rect 13820 18362 13872 18368
rect 13544 18352 13596 18358
rect 13544 18294 13596 18300
rect 13556 17610 13584 18294
rect 13544 17604 13596 17610
rect 13544 17546 13596 17552
rect 13636 17128 13688 17134
rect 13636 17070 13688 17076
rect 13924 17082 13952 19672
rect 14280 19654 14332 19660
rect 14096 19236 14148 19242
rect 14096 19178 14148 19184
rect 14004 18624 14056 18630
rect 14004 18566 14056 18572
rect 14016 18290 14044 18566
rect 14108 18290 14136 19178
rect 14188 18760 14240 18766
rect 14188 18702 14240 18708
rect 14004 18284 14056 18290
rect 14004 18226 14056 18232
rect 14096 18284 14148 18290
rect 14096 18226 14148 18232
rect 14200 17678 14228 18702
rect 14188 17672 14240 17678
rect 14016 17632 14188 17660
rect 14016 17202 14044 17632
rect 14188 17614 14240 17620
rect 14096 17536 14148 17542
rect 14096 17478 14148 17484
rect 14004 17196 14056 17202
rect 14004 17138 14056 17144
rect 13648 16726 13676 17070
rect 13924 17054 14044 17082
rect 13820 16992 13872 16998
rect 13820 16934 13872 16940
rect 13636 16720 13688 16726
rect 13832 16697 13860 16934
rect 13636 16662 13688 16668
rect 13818 16688 13874 16697
rect 13818 16623 13874 16632
rect 13912 16652 13964 16658
rect 13912 16594 13964 16600
rect 13544 16584 13596 16590
rect 13544 16526 13596 16532
rect 13556 16454 13584 16526
rect 13544 16448 13596 16454
rect 13544 16390 13596 16396
rect 13542 16280 13598 16289
rect 13542 16215 13598 16224
rect 13556 16182 13584 16215
rect 13924 16182 13952 16594
rect 14016 16425 14044 17054
rect 14108 16697 14136 17478
rect 14094 16688 14150 16697
rect 14094 16623 14150 16632
rect 14096 16584 14148 16590
rect 14148 16544 14228 16572
rect 14096 16526 14148 16532
rect 14200 16425 14228 16544
rect 14002 16416 14058 16425
rect 14002 16351 14058 16360
rect 14186 16416 14242 16425
rect 14186 16351 14242 16360
rect 13544 16176 13596 16182
rect 13912 16176 13964 16182
rect 13596 16136 13676 16164
rect 13544 16118 13596 16124
rect 13280 16000 13492 16028
rect 12808 15904 12860 15910
rect 12808 15846 12860 15852
rect 12990 15464 13046 15473
rect 12990 15399 13046 15408
rect 12900 14884 12952 14890
rect 12900 14826 12952 14832
rect 12912 14618 12940 14826
rect 12900 14612 12952 14618
rect 12900 14554 12952 14560
rect 12808 13728 12860 13734
rect 12808 13670 12860 13676
rect 12716 12640 12768 12646
rect 12716 12582 12768 12588
rect 12348 12436 12400 12442
rect 12348 12378 12400 12384
rect 11980 12300 12032 12306
rect 11980 12242 12032 12248
rect 11992 11558 12020 12242
rect 12256 11892 12308 11898
rect 12256 11834 12308 11840
rect 12268 11762 12296 11834
rect 12072 11756 12124 11762
rect 12072 11698 12124 11704
rect 12256 11756 12308 11762
rect 12256 11698 12308 11704
rect 11980 11552 12032 11558
rect 11980 11494 12032 11500
rect 11992 10742 12020 11494
rect 12084 11218 12112 11698
rect 12072 11212 12124 11218
rect 12072 11154 12124 11160
rect 12072 11008 12124 11014
rect 12072 10950 12124 10956
rect 11980 10736 12032 10742
rect 11980 10678 12032 10684
rect 12084 9994 12112 10950
rect 12268 10130 12296 11698
rect 12820 11354 12848 13670
rect 12900 13184 12952 13190
rect 12900 13126 12952 13132
rect 12808 11348 12860 11354
rect 12808 11290 12860 11296
rect 12912 11150 12940 13126
rect 13004 11898 13032 15399
rect 13280 14822 13308 16000
rect 13544 15904 13596 15910
rect 13544 15846 13596 15852
rect 13556 15706 13584 15846
rect 13544 15700 13596 15706
rect 13544 15642 13596 15648
rect 13648 15434 13676 16136
rect 13912 16118 13964 16124
rect 14004 16108 14056 16114
rect 14004 16050 14056 16056
rect 14016 15609 14044 16050
rect 14002 15600 14058 15609
rect 14002 15535 14058 15544
rect 13636 15428 13688 15434
rect 13636 15370 13688 15376
rect 14096 15360 14148 15366
rect 14096 15302 14148 15308
rect 13544 15020 13596 15026
rect 13544 14962 13596 14968
rect 13912 15020 13964 15026
rect 13912 14962 13964 14968
rect 13268 14816 13320 14822
rect 13268 14758 13320 14764
rect 13084 14612 13136 14618
rect 13084 14554 13136 14560
rect 13096 14074 13124 14554
rect 13280 14521 13308 14758
rect 13556 14550 13584 14962
rect 13636 14952 13688 14958
rect 13636 14894 13688 14900
rect 13544 14544 13596 14550
rect 13266 14512 13322 14521
rect 13544 14486 13596 14492
rect 13266 14447 13322 14456
rect 13174 14376 13230 14385
rect 13174 14311 13230 14320
rect 13188 14074 13216 14311
rect 13084 14068 13136 14074
rect 13084 14010 13136 14016
rect 13176 14068 13228 14074
rect 13176 14010 13228 14016
rect 13360 13932 13412 13938
rect 13360 13874 13412 13880
rect 13174 13696 13230 13705
rect 13174 13631 13230 13640
rect 13188 13190 13216 13631
rect 13372 13326 13400 13874
rect 13648 13802 13676 14894
rect 13924 14278 13952 14962
rect 13912 14272 13964 14278
rect 13912 14214 13964 14220
rect 13728 13932 13780 13938
rect 13912 13932 13964 13938
rect 13780 13892 13860 13920
rect 13728 13874 13780 13880
rect 13636 13796 13688 13802
rect 13636 13738 13688 13744
rect 13728 13728 13780 13734
rect 13728 13670 13780 13676
rect 13360 13320 13412 13326
rect 13360 13262 13412 13268
rect 13636 13320 13688 13326
rect 13636 13262 13688 13268
rect 13176 13184 13228 13190
rect 13176 13126 13228 13132
rect 13188 12850 13216 13126
rect 13176 12844 13228 12850
rect 13176 12786 13228 12792
rect 13372 12714 13400 13262
rect 13648 12986 13676 13262
rect 13636 12980 13688 12986
rect 13636 12922 13688 12928
rect 13360 12708 13412 12714
rect 13360 12650 13412 12656
rect 13636 12232 13688 12238
rect 13740 12220 13768 13670
rect 13832 13462 13860 13892
rect 13912 13874 13964 13880
rect 13924 13530 13952 13874
rect 13912 13524 13964 13530
rect 13912 13466 13964 13472
rect 13820 13456 13872 13462
rect 13820 13398 13872 13404
rect 14108 12714 14136 15302
rect 14292 15026 14320 19654
rect 14568 19378 14596 20198
rect 14846 20156 15154 20176
rect 14846 20154 14852 20156
rect 14908 20154 14932 20156
rect 14988 20154 15012 20156
rect 15068 20154 15092 20156
rect 15148 20154 15154 20156
rect 14908 20102 14910 20154
rect 15090 20102 15092 20154
rect 14846 20100 14852 20102
rect 14908 20100 14932 20102
rect 14988 20100 15012 20102
rect 15068 20100 15092 20102
rect 15148 20100 15154 20102
rect 14846 20080 15154 20100
rect 15304 19786 15332 20878
rect 15292 19780 15344 19786
rect 15292 19722 15344 19728
rect 14556 19372 14608 19378
rect 14556 19314 14608 19320
rect 14648 19304 14700 19310
rect 14568 19252 14648 19258
rect 14568 19246 14700 19252
rect 14568 19230 14688 19246
rect 14372 18964 14424 18970
rect 14372 18906 14424 18912
rect 14384 18766 14412 18906
rect 14568 18902 14596 19230
rect 14740 19168 14792 19174
rect 14740 19110 14792 19116
rect 15292 19168 15344 19174
rect 15292 19110 15344 19116
rect 14752 18902 14780 19110
rect 14846 19068 15154 19088
rect 14846 19066 14852 19068
rect 14908 19066 14932 19068
rect 14988 19066 15012 19068
rect 15068 19066 15092 19068
rect 15148 19066 15154 19068
rect 14908 19014 14910 19066
rect 15090 19014 15092 19066
rect 14846 19012 14852 19014
rect 14908 19012 14932 19014
rect 14988 19012 15012 19014
rect 15068 19012 15092 19014
rect 15148 19012 15154 19014
rect 14846 18992 15154 19012
rect 14556 18896 14608 18902
rect 14556 18838 14608 18844
rect 14740 18896 14792 18902
rect 14740 18838 14792 18844
rect 14372 18760 14424 18766
rect 14372 18702 14424 18708
rect 14372 18284 14424 18290
rect 14372 18226 14424 18232
rect 14384 16969 14412 18226
rect 14464 18080 14516 18086
rect 14464 18022 14516 18028
rect 14476 17672 14504 18022
rect 14461 17666 14513 17672
rect 14461 17608 14513 17614
rect 14568 17490 14596 18838
rect 15108 18828 15160 18834
rect 15108 18770 15160 18776
rect 14648 18760 14700 18766
rect 14832 18760 14884 18766
rect 14648 18702 14700 18708
rect 14752 18720 14832 18748
rect 14660 18426 14688 18702
rect 14648 18420 14700 18426
rect 14648 18362 14700 18368
rect 14648 17672 14700 17678
rect 14648 17614 14700 17620
rect 14660 17542 14688 17614
rect 14648 17536 14700 17542
rect 14476 17484 14648 17490
rect 14476 17478 14700 17484
rect 14476 17462 14688 17478
rect 14476 17202 14504 17462
rect 14660 17413 14688 17462
rect 14464 17196 14516 17202
rect 14464 17138 14516 17144
rect 14476 17105 14504 17138
rect 14556 17128 14608 17134
rect 14462 17096 14518 17105
rect 14556 17070 14608 17076
rect 14462 17031 14518 17040
rect 14464 16992 14516 16998
rect 14370 16960 14426 16969
rect 14464 16934 14516 16940
rect 14370 16895 14426 16904
rect 14476 16776 14504 16934
rect 14384 16748 14504 16776
rect 14384 16590 14412 16748
rect 14462 16688 14518 16697
rect 14568 16658 14596 17070
rect 14462 16623 14518 16632
rect 14556 16652 14608 16658
rect 14372 16584 14424 16590
rect 14372 16526 14424 16532
rect 14476 16266 14504 16623
rect 14556 16594 14608 16600
rect 14648 16584 14700 16590
rect 14648 16526 14700 16532
rect 14384 16238 14504 16266
rect 14280 15020 14332 15026
rect 14280 14962 14332 14968
rect 14278 14920 14334 14929
rect 14278 14855 14334 14864
rect 14188 14816 14240 14822
rect 14188 14758 14240 14764
rect 14200 14482 14228 14758
rect 14188 14476 14240 14482
rect 14188 14418 14240 14424
rect 14292 14414 14320 14855
rect 14280 14408 14332 14414
rect 14280 14350 14332 14356
rect 14280 14272 14332 14278
rect 14280 14214 14332 14220
rect 14188 13728 14240 13734
rect 14188 13670 14240 13676
rect 14200 13258 14228 13670
rect 14292 13530 14320 14214
rect 14280 13524 14332 13530
rect 14280 13466 14332 13472
rect 14188 13252 14240 13258
rect 14188 13194 14240 13200
rect 14200 12850 14228 13194
rect 14384 12918 14412 16238
rect 14464 16176 14516 16182
rect 14464 16118 14516 16124
rect 14554 16144 14610 16153
rect 14476 15008 14504 16118
rect 14554 16079 14556 16088
rect 14608 16079 14610 16088
rect 14556 16050 14608 16056
rect 14660 15366 14688 16526
rect 14648 15360 14700 15366
rect 14648 15302 14700 15308
rect 14476 14980 14596 15008
rect 14462 14920 14518 14929
rect 14462 14855 14464 14864
rect 14516 14855 14518 14864
rect 14464 14826 14516 14832
rect 14568 14498 14596 14980
rect 14476 14470 14596 14498
rect 14476 14278 14504 14470
rect 14648 14408 14700 14414
rect 14568 14368 14648 14396
rect 14464 14272 14516 14278
rect 14464 14214 14516 14220
rect 14464 13932 14516 13938
rect 14568 13920 14596 14368
rect 14648 14350 14700 14356
rect 14648 14272 14700 14278
rect 14648 14214 14700 14220
rect 14516 13892 14596 13920
rect 14464 13874 14516 13880
rect 14372 12912 14424 12918
rect 14372 12854 14424 12860
rect 14188 12844 14240 12850
rect 14188 12786 14240 12792
rect 14096 12708 14148 12714
rect 14096 12650 14148 12656
rect 14200 12434 14228 12786
rect 14200 12406 14320 12434
rect 13688 12192 13768 12220
rect 13820 12232 13872 12238
rect 13818 12200 13820 12209
rect 13872 12200 13874 12209
rect 13636 12174 13688 12180
rect 12992 11892 13044 11898
rect 12992 11834 13044 11840
rect 12900 11144 12952 11150
rect 12900 11086 12952 11092
rect 13004 11082 13032 11834
rect 13648 11762 13676 12174
rect 13818 12135 13874 12144
rect 13636 11756 13688 11762
rect 13636 11698 13688 11704
rect 13728 11688 13780 11694
rect 13728 11630 13780 11636
rect 13176 11620 13228 11626
rect 13176 11562 13228 11568
rect 13084 11144 13136 11150
rect 13084 11086 13136 11092
rect 12992 11076 13044 11082
rect 12992 11018 13044 11024
rect 12808 10532 12860 10538
rect 12808 10474 12860 10480
rect 12256 10124 12308 10130
rect 12256 10066 12308 10072
rect 12820 10062 12848 10474
rect 12808 10056 12860 10062
rect 12808 9998 12860 10004
rect 12072 9988 12124 9994
rect 12072 9930 12124 9936
rect 11428 9376 11480 9382
rect 11428 9318 11480 9324
rect 11440 9042 11468 9318
rect 11520 9104 11572 9110
rect 11520 9046 11572 9052
rect 11428 9036 11480 9042
rect 11428 8978 11480 8984
rect 11428 8900 11480 8906
rect 11532 8888 11560 9046
rect 11888 9036 11940 9042
rect 11888 8978 11940 8984
rect 11480 8860 11560 8888
rect 11428 8842 11480 8848
rect 11440 8566 11468 8842
rect 11428 8560 11480 8566
rect 11428 8502 11480 8508
rect 11336 6792 11388 6798
rect 11336 6734 11388 6740
rect 11440 6730 11468 8502
rect 11520 8492 11572 8498
rect 11520 8434 11572 8440
rect 11532 8090 11560 8434
rect 11900 8430 11928 8978
rect 11980 8968 12032 8974
rect 11980 8910 12032 8916
rect 11796 8424 11848 8430
rect 11796 8366 11848 8372
rect 11888 8424 11940 8430
rect 11888 8366 11940 8372
rect 11612 8288 11664 8294
rect 11612 8230 11664 8236
rect 11520 8084 11572 8090
rect 11520 8026 11572 8032
rect 11532 7410 11560 8026
rect 11624 7818 11652 8230
rect 11808 7886 11836 8366
rect 11796 7880 11848 7886
rect 11796 7822 11848 7828
rect 11612 7812 11664 7818
rect 11612 7754 11664 7760
rect 11520 7404 11572 7410
rect 11520 7346 11572 7352
rect 11624 7206 11652 7754
rect 11888 7540 11940 7546
rect 11888 7482 11940 7488
rect 11612 7200 11664 7206
rect 11612 7142 11664 7148
rect 11900 6866 11928 7482
rect 11888 6860 11940 6866
rect 11888 6802 11940 6808
rect 11704 6792 11756 6798
rect 11704 6734 11756 6740
rect 11428 6724 11480 6730
rect 11428 6666 11480 6672
rect 11336 6656 11388 6662
rect 11336 6598 11388 6604
rect 11348 5574 11376 6598
rect 11716 5710 11744 6734
rect 11796 6656 11848 6662
rect 11796 6598 11848 6604
rect 11808 5710 11836 6598
rect 11888 6248 11940 6254
rect 11888 6190 11940 6196
rect 11520 5704 11572 5710
rect 11520 5646 11572 5652
rect 11704 5704 11756 5710
rect 11704 5646 11756 5652
rect 11796 5704 11848 5710
rect 11796 5646 11848 5652
rect 11336 5568 11388 5574
rect 11336 5510 11388 5516
rect 11532 5370 11560 5646
rect 11796 5568 11848 5574
rect 11796 5510 11848 5516
rect 11244 5364 11296 5370
rect 11244 5306 11296 5312
rect 11520 5364 11572 5370
rect 11520 5306 11572 5312
rect 11808 5234 11836 5510
rect 11900 5370 11928 6190
rect 11992 6186 12020 8910
rect 12084 8838 12112 9930
rect 12348 9920 12400 9926
rect 12348 9862 12400 9868
rect 12256 9512 12308 9518
rect 12256 9454 12308 9460
rect 12268 8838 12296 9454
rect 12360 9450 12388 9862
rect 13096 9654 13124 11086
rect 13084 9648 13136 9654
rect 13084 9590 13136 9596
rect 12532 9580 12584 9586
rect 12532 9522 12584 9528
rect 12716 9580 12768 9586
rect 12716 9522 12768 9528
rect 12808 9580 12860 9586
rect 12808 9522 12860 9528
rect 12348 9444 12400 9450
rect 12348 9386 12400 9392
rect 12440 9376 12492 9382
rect 12440 9318 12492 9324
rect 12452 8974 12480 9318
rect 12440 8968 12492 8974
rect 12440 8910 12492 8916
rect 12072 8832 12124 8838
rect 12256 8832 12308 8838
rect 12124 8792 12204 8820
rect 12072 8774 12124 8780
rect 12072 8492 12124 8498
rect 12072 8434 12124 8440
rect 12084 8090 12112 8434
rect 12072 8084 12124 8090
rect 12072 8026 12124 8032
rect 12176 7342 12204 8792
rect 12256 8774 12308 8780
rect 12440 8832 12492 8838
rect 12544 8786 12572 9522
rect 12492 8780 12572 8786
rect 12440 8774 12572 8780
rect 12452 8758 12572 8774
rect 12452 8566 12480 8758
rect 12440 8560 12492 8566
rect 12346 8528 12402 8537
rect 12440 8502 12492 8508
rect 12346 8463 12402 8472
rect 12256 8424 12308 8430
rect 12256 8366 12308 8372
rect 12268 7886 12296 8366
rect 12360 8362 12388 8463
rect 12348 8356 12400 8362
rect 12348 8298 12400 8304
rect 12728 8090 12756 9522
rect 12820 8634 12848 9522
rect 13084 8832 13136 8838
rect 13084 8774 13136 8780
rect 12808 8628 12860 8634
rect 12808 8570 12860 8576
rect 12900 8560 12952 8566
rect 12900 8502 12952 8508
rect 12912 8090 12940 8502
rect 13096 8498 13124 8774
rect 13188 8650 13216 11562
rect 13268 11552 13320 11558
rect 13268 11494 13320 11500
rect 13280 11150 13308 11494
rect 13268 11144 13320 11150
rect 13268 11086 13320 11092
rect 13452 11144 13504 11150
rect 13452 11086 13504 11092
rect 13360 11076 13412 11082
rect 13360 11018 13412 11024
rect 13268 10668 13320 10674
rect 13268 10610 13320 10616
rect 13280 10062 13308 10610
rect 13372 10266 13400 11018
rect 13464 10266 13492 11086
rect 13544 10532 13596 10538
rect 13544 10474 13596 10480
rect 13360 10260 13412 10266
rect 13360 10202 13412 10208
rect 13452 10260 13504 10266
rect 13452 10202 13504 10208
rect 13268 10056 13320 10062
rect 13268 9998 13320 10004
rect 13556 8786 13584 10474
rect 13740 9450 13768 11630
rect 13832 11558 13860 12135
rect 14188 12096 14240 12102
rect 14188 12038 14240 12044
rect 14200 11830 14228 12038
rect 14188 11824 14240 11830
rect 14188 11766 14240 11772
rect 13820 11552 13872 11558
rect 13820 11494 13872 11500
rect 13912 11552 13964 11558
rect 13912 11494 13964 11500
rect 13728 9444 13780 9450
rect 13728 9386 13780 9392
rect 13636 9376 13688 9382
rect 13636 9318 13688 9324
rect 13648 9178 13676 9318
rect 13636 9172 13688 9178
rect 13636 9114 13688 9120
rect 13648 8974 13676 9114
rect 13636 8968 13688 8974
rect 13636 8910 13688 8916
rect 13832 8906 13860 11494
rect 13924 11082 13952 11494
rect 14292 11150 14320 12406
rect 14384 11286 14412 12854
rect 14464 12776 14516 12782
rect 14464 12718 14516 12724
rect 14372 11280 14424 11286
rect 14372 11222 14424 11228
rect 14280 11144 14332 11150
rect 14280 11086 14332 11092
rect 13912 11076 13964 11082
rect 13912 11018 13964 11024
rect 13924 10606 13952 11018
rect 14188 10804 14240 10810
rect 14188 10746 14240 10752
rect 13912 10600 13964 10606
rect 13912 10542 13964 10548
rect 13924 9994 13952 10542
rect 14096 10464 14148 10470
rect 14096 10406 14148 10412
rect 13912 9988 13964 9994
rect 13912 9930 13964 9936
rect 14004 9988 14056 9994
rect 14004 9930 14056 9936
rect 14016 9042 14044 9930
rect 14108 9518 14136 10406
rect 14200 10062 14228 10746
rect 14384 10742 14412 11222
rect 14372 10736 14424 10742
rect 14372 10678 14424 10684
rect 14384 10062 14412 10678
rect 14476 10470 14504 12718
rect 14568 12374 14596 13892
rect 14660 13734 14688 14214
rect 14648 13728 14700 13734
rect 14648 13670 14700 13676
rect 14752 13546 14780 18720
rect 14832 18702 14884 18708
rect 15120 18222 15148 18770
rect 15304 18766 15332 19110
rect 15292 18760 15344 18766
rect 15292 18702 15344 18708
rect 15292 18284 15344 18290
rect 15292 18226 15344 18232
rect 15108 18216 15160 18222
rect 15108 18158 15160 18164
rect 14846 17980 15154 18000
rect 14846 17978 14852 17980
rect 14908 17978 14932 17980
rect 14988 17978 15012 17980
rect 15068 17978 15092 17980
rect 15148 17978 15154 17980
rect 14908 17926 14910 17978
rect 15090 17926 15092 17978
rect 14846 17924 14852 17926
rect 14908 17924 14932 17926
rect 14988 17924 15012 17926
rect 15068 17924 15092 17926
rect 15148 17924 15154 17926
rect 14846 17904 15154 17924
rect 15200 17672 15252 17678
rect 15200 17614 15252 17620
rect 15212 16998 15240 17614
rect 15200 16992 15252 16998
rect 15200 16934 15252 16940
rect 14846 16892 15154 16912
rect 14846 16890 14852 16892
rect 14908 16890 14932 16892
rect 14988 16890 15012 16892
rect 15068 16890 15092 16892
rect 15148 16890 15154 16892
rect 14908 16838 14910 16890
rect 15090 16838 15092 16890
rect 14846 16836 14852 16838
rect 14908 16836 14932 16838
rect 14988 16836 15012 16838
rect 15068 16836 15092 16838
rect 15148 16836 15154 16838
rect 14846 16816 15154 16836
rect 15016 16720 15068 16726
rect 15016 16662 15068 16668
rect 15028 15978 15056 16662
rect 15108 16584 15160 16590
rect 15160 16544 15240 16572
rect 15108 16526 15160 16532
rect 15212 16454 15240 16544
rect 15108 16448 15160 16454
rect 15200 16448 15252 16454
rect 15108 16390 15160 16396
rect 15198 16416 15200 16425
rect 15252 16416 15254 16425
rect 15120 16114 15148 16390
rect 15198 16351 15254 16360
rect 15108 16108 15160 16114
rect 15108 16050 15160 16056
rect 15200 16108 15252 16114
rect 15200 16050 15252 16056
rect 15016 15972 15068 15978
rect 15016 15914 15068 15920
rect 14846 15804 15154 15824
rect 14846 15802 14852 15804
rect 14908 15802 14932 15804
rect 14988 15802 15012 15804
rect 15068 15802 15092 15804
rect 15148 15802 15154 15804
rect 14908 15750 14910 15802
rect 15090 15750 15092 15802
rect 14846 15748 14852 15750
rect 14908 15748 14932 15750
rect 14988 15748 15012 15750
rect 15068 15748 15092 15750
rect 15148 15748 15154 15750
rect 14846 15728 15154 15748
rect 15212 15706 15240 16050
rect 15200 15700 15252 15706
rect 15200 15642 15252 15648
rect 15016 15428 15068 15434
rect 15016 15370 15068 15376
rect 15028 15162 15056 15370
rect 15016 15156 15068 15162
rect 15016 15098 15068 15104
rect 15200 15020 15252 15026
rect 15200 14962 15252 14968
rect 14846 14716 15154 14736
rect 14846 14714 14852 14716
rect 14908 14714 14932 14716
rect 14988 14714 15012 14716
rect 15068 14714 15092 14716
rect 15148 14714 15154 14716
rect 14908 14662 14910 14714
rect 15090 14662 15092 14714
rect 14846 14660 14852 14662
rect 14908 14660 14932 14662
rect 14988 14660 15012 14662
rect 15068 14660 15092 14662
rect 15148 14660 15154 14662
rect 14846 14640 15154 14660
rect 15212 14521 15240 14962
rect 15198 14512 15254 14521
rect 15198 14447 15254 14456
rect 15200 14340 15252 14346
rect 15200 14282 15252 14288
rect 15212 14074 15240 14282
rect 15200 14068 15252 14074
rect 15200 14010 15252 14016
rect 14846 13628 15154 13648
rect 14846 13626 14852 13628
rect 14908 13626 14932 13628
rect 14988 13626 15012 13628
rect 15068 13626 15092 13628
rect 15148 13626 15154 13628
rect 14908 13574 14910 13626
rect 15090 13574 15092 13626
rect 14846 13572 14852 13574
rect 14908 13572 14932 13574
rect 14988 13572 15012 13574
rect 15068 13572 15092 13574
rect 15148 13572 15154 13574
rect 14846 13552 15154 13572
rect 14660 13518 14780 13546
rect 15200 13524 15252 13530
rect 14660 12782 14688 13518
rect 15200 13466 15252 13472
rect 14740 13456 14792 13462
rect 14740 13398 14792 13404
rect 14648 12776 14700 12782
rect 14648 12718 14700 12724
rect 14648 12640 14700 12646
rect 14648 12582 14700 12588
rect 14556 12368 14608 12374
rect 14556 12310 14608 12316
rect 14660 12238 14688 12582
rect 14752 12345 14780 13398
rect 14846 12540 15154 12560
rect 14846 12538 14852 12540
rect 14908 12538 14932 12540
rect 14988 12538 15012 12540
rect 15068 12538 15092 12540
rect 15148 12538 15154 12540
rect 14908 12486 14910 12538
rect 15090 12486 15092 12538
rect 14846 12484 14852 12486
rect 14908 12484 14932 12486
rect 14988 12484 15012 12486
rect 15068 12484 15092 12486
rect 15148 12484 15154 12486
rect 14846 12464 15154 12484
rect 14832 12368 14884 12374
rect 14738 12336 14794 12345
rect 14832 12310 14884 12316
rect 14738 12271 14794 12280
rect 14844 12238 14872 12310
rect 15212 12306 15240 13466
rect 15304 12850 15332 18226
rect 15396 16561 15424 22066
rect 15764 21486 15792 22066
rect 15856 22066 15976 22094
rect 16304 22092 16356 22098
rect 15856 21554 15884 22066
rect 16304 22034 16356 22040
rect 15844 21548 15896 21554
rect 15844 21490 15896 21496
rect 15752 21480 15804 21486
rect 15752 21422 15804 21428
rect 15568 21344 15620 21350
rect 15568 21286 15620 21292
rect 15476 20596 15528 20602
rect 15476 20538 15528 20544
rect 15488 20058 15516 20538
rect 15580 20466 15608 21286
rect 15764 21146 15792 21422
rect 15752 21140 15804 21146
rect 15752 21082 15804 21088
rect 16316 21010 16344 22034
rect 16488 21956 16540 21962
rect 16488 21898 16540 21904
rect 16500 21690 16528 21898
rect 16684 21894 16712 22170
rect 17052 21894 17080 22918
rect 17144 22710 17172 22918
rect 17224 22772 17276 22778
rect 17224 22714 17276 22720
rect 17132 22704 17184 22710
rect 17132 22646 17184 22652
rect 17144 22030 17172 22646
rect 17236 22030 17264 22714
rect 17972 22642 18000 22918
rect 17960 22636 18012 22642
rect 17960 22578 18012 22584
rect 17592 22228 17644 22234
rect 17592 22170 17644 22176
rect 17604 22030 17632 22170
rect 17132 22024 17184 22030
rect 17132 21966 17184 21972
rect 17224 22024 17276 22030
rect 17224 21966 17276 21972
rect 17592 22024 17644 22030
rect 17592 21966 17644 21972
rect 16580 21888 16632 21894
rect 16580 21830 16632 21836
rect 16672 21888 16724 21894
rect 16672 21830 16724 21836
rect 17040 21888 17092 21894
rect 17040 21830 17092 21836
rect 16488 21684 16540 21690
rect 16488 21626 16540 21632
rect 16592 21350 16620 21830
rect 16580 21344 16632 21350
rect 16580 21286 16632 21292
rect 16304 21004 16356 21010
rect 16304 20946 16356 20952
rect 16120 20800 16172 20806
rect 16120 20742 16172 20748
rect 15568 20460 15620 20466
rect 15568 20402 15620 20408
rect 15476 20052 15528 20058
rect 15476 19994 15528 20000
rect 15488 19514 15516 19994
rect 15476 19508 15528 19514
rect 15476 19450 15528 19456
rect 15476 18216 15528 18222
rect 15476 18158 15528 18164
rect 15488 17746 15516 18158
rect 15476 17740 15528 17746
rect 15476 17682 15528 17688
rect 15488 17134 15516 17682
rect 15580 17338 15608 20402
rect 16132 20262 16160 20742
rect 16316 20534 16344 20946
rect 16304 20528 16356 20534
rect 16304 20470 16356 20476
rect 16120 20256 16172 20262
rect 16120 20198 16172 20204
rect 16132 19854 16160 20198
rect 16212 20052 16264 20058
rect 16212 19994 16264 20000
rect 16120 19848 16172 19854
rect 16120 19790 16172 19796
rect 16028 19780 16080 19786
rect 16028 19722 16080 19728
rect 15752 19712 15804 19718
rect 15752 19654 15804 19660
rect 15660 18624 15712 18630
rect 15660 18566 15712 18572
rect 15672 17678 15700 18566
rect 15764 18358 15792 19654
rect 16040 19378 16068 19722
rect 16224 19514 16252 19994
rect 16580 19848 16632 19854
rect 16580 19790 16632 19796
rect 16212 19508 16264 19514
rect 16212 19450 16264 19456
rect 16592 19378 16620 19790
rect 16028 19372 16080 19378
rect 16028 19314 16080 19320
rect 16580 19372 16632 19378
rect 16580 19314 16632 19320
rect 15936 19168 15988 19174
rect 15936 19110 15988 19116
rect 15752 18352 15804 18358
rect 15752 18294 15804 18300
rect 15660 17672 15712 17678
rect 15660 17614 15712 17620
rect 15568 17332 15620 17338
rect 15568 17274 15620 17280
rect 15752 17196 15804 17202
rect 15752 17138 15804 17144
rect 15476 17128 15528 17134
rect 15476 17070 15528 17076
rect 15764 16658 15792 17138
rect 15844 16788 15896 16794
rect 15844 16730 15896 16736
rect 15752 16652 15804 16658
rect 15752 16594 15804 16600
rect 15476 16584 15528 16590
rect 15382 16552 15438 16561
rect 15476 16526 15528 16532
rect 15660 16584 15712 16590
rect 15660 16526 15712 16532
rect 15382 16487 15438 16496
rect 15488 16250 15516 16526
rect 15476 16244 15528 16250
rect 15476 16186 15528 16192
rect 15382 16008 15438 16017
rect 15382 15943 15384 15952
rect 15436 15943 15438 15952
rect 15384 15914 15436 15920
rect 15382 15600 15438 15609
rect 15382 15535 15438 15544
rect 15396 15366 15424 15535
rect 15384 15360 15436 15366
rect 15384 15302 15436 15308
rect 15396 14414 15424 15302
rect 15568 15088 15620 15094
rect 15568 15030 15620 15036
rect 15476 15020 15528 15026
rect 15476 14962 15528 14968
rect 15488 14618 15516 14962
rect 15580 14618 15608 15030
rect 15476 14612 15528 14618
rect 15476 14554 15528 14560
rect 15568 14612 15620 14618
rect 15568 14554 15620 14560
rect 15476 14476 15528 14482
rect 15476 14418 15528 14424
rect 15384 14408 15436 14414
rect 15384 14350 15436 14356
rect 15384 14068 15436 14074
rect 15384 14010 15436 14016
rect 15292 12844 15344 12850
rect 15292 12786 15344 12792
rect 15396 12442 15424 14010
rect 15384 12436 15436 12442
rect 15384 12378 15436 12384
rect 15200 12300 15252 12306
rect 15200 12242 15252 12248
rect 14648 12232 14700 12238
rect 14648 12174 14700 12180
rect 14832 12232 14884 12238
rect 14832 12174 14884 12180
rect 15212 11937 15240 12242
rect 15198 11928 15254 11937
rect 15198 11863 15254 11872
rect 14846 11452 15154 11472
rect 14846 11450 14852 11452
rect 14908 11450 14932 11452
rect 14988 11450 15012 11452
rect 15068 11450 15092 11452
rect 15148 11450 15154 11452
rect 14908 11398 14910 11450
rect 15090 11398 15092 11450
rect 14846 11396 14852 11398
rect 14908 11396 14932 11398
rect 14988 11396 15012 11398
rect 15068 11396 15092 11398
rect 15148 11396 15154 11398
rect 14846 11376 15154 11396
rect 14556 11280 14608 11286
rect 14556 11222 14608 11228
rect 15014 11248 15070 11257
rect 14464 10464 14516 10470
rect 14464 10406 14516 10412
rect 14188 10056 14240 10062
rect 14188 9998 14240 10004
rect 14372 10056 14424 10062
rect 14372 9998 14424 10004
rect 14096 9512 14148 9518
rect 14096 9454 14148 9460
rect 14004 9036 14056 9042
rect 14004 8978 14056 8984
rect 13820 8900 13872 8906
rect 13820 8842 13872 8848
rect 13556 8758 13676 8786
rect 13188 8622 13400 8650
rect 13084 8492 13136 8498
rect 13084 8434 13136 8440
rect 13268 8492 13320 8498
rect 13268 8434 13320 8440
rect 12716 8084 12768 8090
rect 12716 8026 12768 8032
rect 12900 8084 12952 8090
rect 12900 8026 12952 8032
rect 13096 7954 13124 8434
rect 13176 8288 13228 8294
rect 13176 8230 13228 8236
rect 12440 7948 12492 7954
rect 12440 7890 12492 7896
rect 13084 7948 13136 7954
rect 13084 7890 13136 7896
rect 12256 7880 12308 7886
rect 12256 7822 12308 7828
rect 12452 7410 12480 7890
rect 12440 7404 12492 7410
rect 12440 7346 12492 7352
rect 12624 7404 12676 7410
rect 12624 7346 12676 7352
rect 12164 7336 12216 7342
rect 12636 7290 12664 7346
rect 13188 7342 13216 8230
rect 13280 7886 13308 8434
rect 13372 7954 13400 8622
rect 13360 7948 13412 7954
rect 13360 7890 13412 7896
rect 13268 7880 13320 7886
rect 13268 7822 13320 7828
rect 13280 7478 13308 7822
rect 13648 7818 13676 8758
rect 14016 8498 14044 8978
rect 14004 8492 14056 8498
rect 14004 8434 14056 8440
rect 14108 8430 14136 9454
rect 14096 8424 14148 8430
rect 14096 8366 14148 8372
rect 14108 8072 14136 8366
rect 14200 8294 14228 9998
rect 14280 9920 14332 9926
rect 14280 9862 14332 9868
rect 14292 8498 14320 9862
rect 14476 9586 14504 10406
rect 14464 9580 14516 9586
rect 14464 9522 14516 9528
rect 14464 8900 14516 8906
rect 14464 8842 14516 8848
rect 14476 8498 14504 8842
rect 14280 8492 14332 8498
rect 14464 8492 14516 8498
rect 14280 8434 14332 8440
rect 14384 8452 14464 8480
rect 14188 8288 14240 8294
rect 14188 8230 14240 8236
rect 14188 8084 14240 8090
rect 14108 8044 14188 8072
rect 14188 8026 14240 8032
rect 14292 7818 14320 8434
rect 13636 7812 13688 7818
rect 13636 7754 13688 7760
rect 14280 7812 14332 7818
rect 14280 7754 14332 7760
rect 13268 7472 13320 7478
rect 13268 7414 13320 7420
rect 12164 7278 12216 7284
rect 12544 7262 12664 7290
rect 13176 7336 13228 7342
rect 13176 7278 13228 7284
rect 12900 7268 12952 7274
rect 12544 7002 12572 7262
rect 12900 7210 12952 7216
rect 12532 6996 12584 7002
rect 12532 6938 12584 6944
rect 12164 6928 12216 6934
rect 12164 6870 12216 6876
rect 11980 6180 12032 6186
rect 11980 6122 12032 6128
rect 11888 5364 11940 5370
rect 11888 5306 11940 5312
rect 11796 5228 11848 5234
rect 11796 5170 11848 5176
rect 11060 5024 11112 5030
rect 11060 4966 11112 4972
rect 11704 5024 11756 5030
rect 11704 4966 11756 4972
rect 11612 4684 11664 4690
rect 11612 4626 11664 4632
rect 11428 4616 11480 4622
rect 11428 4558 11480 4564
rect 11440 4010 11468 4558
rect 11428 4004 11480 4010
rect 11428 3946 11480 3952
rect 10876 3528 10928 3534
rect 8206 3496 8262 3505
rect 10876 3470 10928 3476
rect 11440 3466 11468 3946
rect 11624 3942 11652 4626
rect 11716 4282 11744 4966
rect 11704 4276 11756 4282
rect 11704 4218 11756 4224
rect 11612 3936 11664 3942
rect 11612 3878 11664 3884
rect 11796 3936 11848 3942
rect 11796 3878 11848 3884
rect 11624 3466 11652 3878
rect 11808 3534 11836 3878
rect 11900 3534 11928 5306
rect 11796 3528 11848 3534
rect 11796 3470 11848 3476
rect 11888 3528 11940 3534
rect 11888 3470 11940 3476
rect 8206 3431 8262 3440
rect 11428 3460 11480 3466
rect 8220 3194 8248 3431
rect 11428 3402 11480 3408
rect 11612 3460 11664 3466
rect 11612 3402 11664 3408
rect 10968 3392 11020 3398
rect 10968 3334 11020 3340
rect 10214 3292 10522 3312
rect 10214 3290 10220 3292
rect 10276 3290 10300 3292
rect 10356 3290 10380 3292
rect 10436 3290 10460 3292
rect 10516 3290 10522 3292
rect 10276 3238 10278 3290
rect 10458 3238 10460 3290
rect 10214 3236 10220 3238
rect 10276 3236 10300 3238
rect 10356 3236 10380 3238
rect 10436 3236 10460 3238
rect 10516 3236 10522 3238
rect 10214 3216 10522 3236
rect 8208 3188 8260 3194
rect 8208 3130 8260 3136
rect 8116 3052 8168 3058
rect 8116 2994 8168 3000
rect 10980 2990 11008 3334
rect 11992 3194 12020 6122
rect 12072 6112 12124 6118
rect 12072 6054 12124 6060
rect 12084 5710 12112 6054
rect 12072 5704 12124 5710
rect 12072 5646 12124 5652
rect 12176 5642 12204 6870
rect 12440 6656 12492 6662
rect 12440 6598 12492 6604
rect 12256 6316 12308 6322
rect 12256 6258 12308 6264
rect 12268 5914 12296 6258
rect 12348 6112 12400 6118
rect 12348 6054 12400 6060
rect 12256 5908 12308 5914
rect 12256 5850 12308 5856
rect 12360 5846 12388 6054
rect 12348 5840 12400 5846
rect 12348 5782 12400 5788
rect 12452 5710 12480 6598
rect 12544 5846 12572 6938
rect 12912 6798 12940 7210
rect 12716 6792 12768 6798
rect 12716 6734 12768 6740
rect 12900 6792 12952 6798
rect 12900 6734 12952 6740
rect 12728 6458 12756 6734
rect 12808 6656 12860 6662
rect 12808 6598 12860 6604
rect 12716 6452 12768 6458
rect 12636 6412 12716 6440
rect 12532 5840 12584 5846
rect 12532 5782 12584 5788
rect 12440 5704 12492 5710
rect 12440 5646 12492 5652
rect 12164 5636 12216 5642
rect 12164 5578 12216 5584
rect 12176 5234 12204 5578
rect 12256 5296 12308 5302
rect 12256 5238 12308 5244
rect 12164 5228 12216 5234
rect 12164 5170 12216 5176
rect 12176 4622 12204 5170
rect 12268 5137 12296 5238
rect 12254 5128 12310 5137
rect 12254 5063 12310 5072
rect 12452 5030 12480 5646
rect 12636 5166 12664 6412
rect 12716 6394 12768 6400
rect 12716 5840 12768 5846
rect 12716 5782 12768 5788
rect 12624 5160 12676 5166
rect 12624 5102 12676 5108
rect 12440 5024 12492 5030
rect 12440 4966 12492 4972
rect 12530 4992 12586 5001
rect 12530 4927 12586 4936
rect 12256 4752 12308 4758
rect 12256 4694 12308 4700
rect 12164 4616 12216 4622
rect 12164 4558 12216 4564
rect 12268 4146 12296 4694
rect 12164 4140 12216 4146
rect 12164 4082 12216 4088
rect 12256 4140 12308 4146
rect 12256 4082 12308 4088
rect 12176 3942 12204 4082
rect 12164 3936 12216 3942
rect 12164 3878 12216 3884
rect 12256 3664 12308 3670
rect 12544 3618 12572 4927
rect 12636 4826 12664 5102
rect 12624 4820 12676 4826
rect 12624 4762 12676 4768
rect 12728 4706 12756 5782
rect 12636 4678 12756 4706
rect 12636 4622 12664 4678
rect 12624 4616 12676 4622
rect 12624 4558 12676 4564
rect 12624 4480 12676 4486
rect 12624 4422 12676 4428
rect 12636 4146 12664 4422
rect 12820 4282 12848 6598
rect 12900 5908 12952 5914
rect 12900 5850 12952 5856
rect 12912 5234 12940 5850
rect 13188 5778 13216 7278
rect 13648 6798 13676 7754
rect 14384 7410 14412 8452
rect 14464 8434 14516 8440
rect 14464 8288 14516 8294
rect 14464 8230 14516 8236
rect 14476 7546 14504 8230
rect 14464 7540 14516 7546
rect 14464 7482 14516 7488
rect 14372 7404 14424 7410
rect 14372 7346 14424 7352
rect 14372 7200 14424 7206
rect 14372 7142 14424 7148
rect 13636 6792 13688 6798
rect 13636 6734 13688 6740
rect 13912 6792 13964 6798
rect 13912 6734 13964 6740
rect 13924 6390 13952 6734
rect 14188 6724 14240 6730
rect 14188 6666 14240 6672
rect 14004 6656 14056 6662
rect 14004 6598 14056 6604
rect 13912 6384 13964 6390
rect 13912 6326 13964 6332
rect 14016 6322 14044 6598
rect 14200 6458 14228 6666
rect 14188 6452 14240 6458
rect 14188 6394 14240 6400
rect 14384 6322 14412 7142
rect 14004 6316 14056 6322
rect 14004 6258 14056 6264
rect 14372 6316 14424 6322
rect 14372 6258 14424 6264
rect 13360 5908 13412 5914
rect 13360 5850 13412 5856
rect 13176 5772 13228 5778
rect 13176 5714 13228 5720
rect 13084 5636 13136 5642
rect 13084 5578 13136 5584
rect 12900 5228 12952 5234
rect 12900 5170 12952 5176
rect 13096 5166 13124 5578
rect 13084 5160 13136 5166
rect 13084 5102 13136 5108
rect 12900 5024 12952 5030
rect 12900 4966 12952 4972
rect 12912 4690 12940 4966
rect 12992 4820 13044 4826
rect 12992 4762 13044 4768
rect 12900 4684 12952 4690
rect 12900 4626 12952 4632
rect 12808 4276 12860 4282
rect 12808 4218 12860 4224
rect 12624 4140 12676 4146
rect 12624 4082 12676 4088
rect 12900 4140 12952 4146
rect 12900 4082 12952 4088
rect 12308 3612 12572 3618
rect 12256 3606 12572 3612
rect 12268 3596 12572 3606
rect 12268 3590 12440 3596
rect 12492 3590 12572 3596
rect 12440 3538 12492 3544
rect 12636 3534 12664 4082
rect 12912 3942 12940 4082
rect 13004 4078 13032 4762
rect 12992 4072 13044 4078
rect 12992 4014 13044 4020
rect 12900 3936 12952 3942
rect 12900 3878 12952 3884
rect 13096 3738 13124 5102
rect 13188 5030 13216 5714
rect 13372 5642 13400 5850
rect 13912 5704 13964 5710
rect 13912 5646 13964 5652
rect 13360 5636 13412 5642
rect 13360 5578 13412 5584
rect 13360 5228 13412 5234
rect 13360 5170 13412 5176
rect 13176 5024 13228 5030
rect 13176 4966 13228 4972
rect 13372 4758 13400 5170
rect 13924 5166 13952 5646
rect 14016 5234 14044 6258
rect 14568 5642 14596 11222
rect 15212 11218 15240 11863
rect 15292 11756 15344 11762
rect 15292 11698 15344 11704
rect 15014 11183 15016 11192
rect 15068 11183 15070 11192
rect 15200 11212 15252 11218
rect 15016 11154 15068 11160
rect 15200 11154 15252 11160
rect 14648 11144 14700 11150
rect 14648 11086 14700 11092
rect 14660 9994 14688 11086
rect 15200 11076 15252 11082
rect 15200 11018 15252 11024
rect 15212 10470 15240 11018
rect 15304 10674 15332 11698
rect 15488 11354 15516 14418
rect 15580 13530 15608 14554
rect 15672 14550 15700 16526
rect 15764 16046 15792 16594
rect 15752 16040 15804 16046
rect 15752 15982 15804 15988
rect 15856 15502 15884 16730
rect 15948 16590 15976 19110
rect 16040 18766 16068 19314
rect 16592 18766 16620 19314
rect 16028 18760 16080 18766
rect 16028 18702 16080 18708
rect 16580 18760 16632 18766
rect 16580 18702 16632 18708
rect 16040 18290 16068 18702
rect 16684 18698 16712 21830
rect 16764 21072 16816 21078
rect 16764 21014 16816 21020
rect 16776 20466 16804 21014
rect 16764 20460 16816 20466
rect 16764 20402 16816 20408
rect 17052 19514 17080 21830
rect 17144 21554 17172 21966
rect 17960 21888 18012 21894
rect 17960 21830 18012 21836
rect 17132 21548 17184 21554
rect 17132 21490 17184 21496
rect 17144 20534 17172 21490
rect 17224 21344 17276 21350
rect 17222 21312 17224 21321
rect 17276 21312 17278 21321
rect 17222 21247 17278 21256
rect 17132 20528 17184 20534
rect 17132 20470 17184 20476
rect 17972 19854 18000 21830
rect 18248 21622 18276 22918
rect 18236 21616 18288 21622
rect 18236 21558 18288 21564
rect 18340 20602 18368 27406
rect 25044 27396 25096 27402
rect 25044 27338 25096 27344
rect 22836 27328 22888 27334
rect 22836 27270 22888 27276
rect 23480 27328 23532 27334
rect 23480 27270 23532 27276
rect 19478 27228 19786 27248
rect 19478 27226 19484 27228
rect 19540 27226 19564 27228
rect 19620 27226 19644 27228
rect 19700 27226 19724 27228
rect 19780 27226 19786 27228
rect 19540 27174 19542 27226
rect 19722 27174 19724 27226
rect 19478 27172 19484 27174
rect 19540 27172 19564 27174
rect 19620 27172 19644 27174
rect 19700 27172 19724 27174
rect 19780 27172 19786 27174
rect 19478 27152 19786 27172
rect 22376 26988 22428 26994
rect 22376 26930 22428 26936
rect 20904 26920 20956 26926
rect 20904 26862 20956 26868
rect 19478 26140 19786 26160
rect 19478 26138 19484 26140
rect 19540 26138 19564 26140
rect 19620 26138 19644 26140
rect 19700 26138 19724 26140
rect 19780 26138 19786 26140
rect 19540 26086 19542 26138
rect 19722 26086 19724 26138
rect 19478 26084 19484 26086
rect 19540 26084 19564 26086
rect 19620 26084 19644 26086
rect 19700 26084 19724 26086
rect 19780 26084 19786 26086
rect 19478 26064 19786 26084
rect 19478 25052 19786 25072
rect 19478 25050 19484 25052
rect 19540 25050 19564 25052
rect 19620 25050 19644 25052
rect 19700 25050 19724 25052
rect 19780 25050 19786 25052
rect 19540 24998 19542 25050
rect 19722 24998 19724 25050
rect 19478 24996 19484 24998
rect 19540 24996 19564 24998
rect 19620 24996 19644 24998
rect 19700 24996 19724 24998
rect 19780 24996 19786 24998
rect 19478 24976 19786 24996
rect 19478 23964 19786 23984
rect 19478 23962 19484 23964
rect 19540 23962 19564 23964
rect 19620 23962 19644 23964
rect 19700 23962 19724 23964
rect 19780 23962 19786 23964
rect 19540 23910 19542 23962
rect 19722 23910 19724 23962
rect 19478 23908 19484 23910
rect 19540 23908 19564 23910
rect 19620 23908 19644 23910
rect 19700 23908 19724 23910
rect 19780 23908 19786 23910
rect 19478 23888 19786 23908
rect 20916 23798 20944 26862
rect 20904 23792 20956 23798
rect 20904 23734 20956 23740
rect 19248 23588 19300 23594
rect 19248 23530 19300 23536
rect 18420 23112 18472 23118
rect 18420 23054 18472 23060
rect 18880 23112 18932 23118
rect 18880 23054 18932 23060
rect 18432 21690 18460 23054
rect 18696 22976 18748 22982
rect 18696 22918 18748 22924
rect 18708 22710 18736 22918
rect 18696 22704 18748 22710
rect 18696 22646 18748 22652
rect 18892 22234 18920 23054
rect 19260 23050 19288 23530
rect 20536 23316 20588 23322
rect 20536 23258 20588 23264
rect 19984 23112 20036 23118
rect 19984 23054 20036 23060
rect 20260 23112 20312 23118
rect 20260 23054 20312 23060
rect 19248 23044 19300 23050
rect 19248 22986 19300 22992
rect 19340 23044 19392 23050
rect 19340 22986 19392 22992
rect 19892 23044 19944 23050
rect 19892 22986 19944 22992
rect 19352 22642 19380 22986
rect 19478 22876 19786 22896
rect 19478 22874 19484 22876
rect 19540 22874 19564 22876
rect 19620 22874 19644 22876
rect 19700 22874 19724 22876
rect 19780 22874 19786 22876
rect 19540 22822 19542 22874
rect 19722 22822 19724 22874
rect 19478 22820 19484 22822
rect 19540 22820 19564 22822
rect 19620 22820 19644 22822
rect 19700 22820 19724 22822
rect 19780 22820 19786 22822
rect 19478 22800 19786 22820
rect 19340 22636 19392 22642
rect 19340 22578 19392 22584
rect 19064 22432 19116 22438
rect 19064 22374 19116 22380
rect 19708 22432 19760 22438
rect 19708 22374 19760 22380
rect 18880 22228 18932 22234
rect 18880 22170 18932 22176
rect 19076 22166 19104 22374
rect 18788 22160 18840 22166
rect 18788 22102 18840 22108
rect 19064 22160 19116 22166
rect 19064 22102 19116 22108
rect 18604 22024 18656 22030
rect 18604 21966 18656 21972
rect 18696 22024 18748 22030
rect 18696 21966 18748 21972
rect 18420 21684 18472 21690
rect 18420 21626 18472 21632
rect 18616 21622 18644 21966
rect 18708 21894 18736 21966
rect 18800 21962 18828 22102
rect 18972 22092 19024 22098
rect 18972 22034 19024 22040
rect 18984 21978 19012 22034
rect 19076 21978 19104 22102
rect 18788 21956 18840 21962
rect 18984 21950 19104 21978
rect 19720 21962 19748 22374
rect 19904 22098 19932 22986
rect 19892 22092 19944 22098
rect 19892 22034 19944 22040
rect 19904 21962 19932 22034
rect 19708 21956 19760 21962
rect 18788 21898 18840 21904
rect 19708 21898 19760 21904
rect 19892 21956 19944 21962
rect 19892 21898 19944 21904
rect 18696 21888 18748 21894
rect 18696 21830 18748 21836
rect 19340 21888 19392 21894
rect 19340 21830 19392 21836
rect 18604 21616 18656 21622
rect 18604 21558 18656 21564
rect 18880 21548 18932 21554
rect 18880 21490 18932 21496
rect 18420 21344 18472 21350
rect 18420 21286 18472 21292
rect 18432 21010 18460 21286
rect 18892 21146 18920 21490
rect 19352 21321 19380 21830
rect 19478 21788 19786 21808
rect 19478 21786 19484 21788
rect 19540 21786 19564 21788
rect 19620 21786 19644 21788
rect 19700 21786 19724 21788
rect 19780 21786 19786 21788
rect 19540 21734 19542 21786
rect 19722 21734 19724 21786
rect 19478 21732 19484 21734
rect 19540 21732 19564 21734
rect 19620 21732 19644 21734
rect 19700 21732 19724 21734
rect 19780 21732 19786 21734
rect 19478 21712 19786 21732
rect 19616 21548 19668 21554
rect 19616 21490 19668 21496
rect 19338 21312 19394 21321
rect 19338 21247 19394 21256
rect 18880 21140 18932 21146
rect 18880 21082 18932 21088
rect 19628 21010 19656 21490
rect 18420 21004 18472 21010
rect 18420 20946 18472 20952
rect 19340 21004 19392 21010
rect 19340 20946 19392 20952
rect 19616 21004 19668 21010
rect 19616 20946 19668 20952
rect 18328 20596 18380 20602
rect 18328 20538 18380 20544
rect 18432 20482 18460 20946
rect 19248 20800 19300 20806
rect 19248 20742 19300 20748
rect 18340 20454 18460 20482
rect 18788 20460 18840 20466
rect 18340 19854 18368 20454
rect 18788 20402 18840 20408
rect 19156 20460 19208 20466
rect 19156 20402 19208 20408
rect 18420 20256 18472 20262
rect 18420 20198 18472 20204
rect 18432 19854 18460 20198
rect 17684 19848 17736 19854
rect 17684 19790 17736 19796
rect 17960 19848 18012 19854
rect 17960 19790 18012 19796
rect 18328 19848 18380 19854
rect 18328 19790 18380 19796
rect 18420 19848 18472 19854
rect 18420 19790 18472 19796
rect 17408 19712 17460 19718
rect 17408 19654 17460 19660
rect 17040 19508 17092 19514
rect 17040 19450 17092 19456
rect 16764 19168 16816 19174
rect 16764 19110 16816 19116
rect 16776 18970 16804 19110
rect 16764 18964 16816 18970
rect 16764 18906 16816 18912
rect 17316 18828 17368 18834
rect 17316 18770 17368 18776
rect 16948 18760 17000 18766
rect 16948 18702 17000 18708
rect 16672 18692 16724 18698
rect 16672 18634 16724 18640
rect 16212 18624 16264 18630
rect 16212 18566 16264 18572
rect 16028 18284 16080 18290
rect 16028 18226 16080 18232
rect 16120 17536 16172 17542
rect 16120 17478 16172 17484
rect 16132 17202 16160 17478
rect 16120 17196 16172 17202
rect 16120 17138 16172 17144
rect 15936 16584 15988 16590
rect 15936 16526 15988 16532
rect 16028 16108 16080 16114
rect 16028 16050 16080 16056
rect 16040 15502 16068 16050
rect 16120 16040 16172 16046
rect 16120 15982 16172 15988
rect 15844 15496 15896 15502
rect 15844 15438 15896 15444
rect 16028 15496 16080 15502
rect 16028 15438 16080 15444
rect 16040 15094 16068 15438
rect 16028 15088 16080 15094
rect 16028 15030 16080 15036
rect 15752 14952 15804 14958
rect 15752 14894 15804 14900
rect 15660 14544 15712 14550
rect 15660 14486 15712 14492
rect 15764 14396 15792 14894
rect 15844 14884 15896 14890
rect 15844 14826 15896 14832
rect 15672 14368 15792 14396
rect 15672 13938 15700 14368
rect 15752 14272 15804 14278
rect 15752 14214 15804 14220
rect 15660 13932 15712 13938
rect 15660 13874 15712 13880
rect 15568 13524 15620 13530
rect 15568 13466 15620 13472
rect 15568 13320 15620 13326
rect 15672 13308 15700 13874
rect 15764 13326 15792 14214
rect 15856 14006 15884 14826
rect 16040 14482 16068 15030
rect 16132 14482 16160 15982
rect 16224 15162 16252 18566
rect 16960 18290 16988 18702
rect 17328 18358 17356 18770
rect 17420 18766 17448 19654
rect 17696 18766 17724 19790
rect 18236 19780 18288 19786
rect 18236 19722 18288 19728
rect 17776 19372 17828 19378
rect 17776 19314 17828 19320
rect 17788 18970 17816 19314
rect 17776 18964 17828 18970
rect 17776 18906 17828 18912
rect 17776 18828 17828 18834
rect 17776 18770 17828 18776
rect 17408 18760 17460 18766
rect 17408 18702 17460 18708
rect 17684 18760 17736 18766
rect 17684 18702 17736 18708
rect 17040 18352 17092 18358
rect 17040 18294 17092 18300
rect 17316 18352 17368 18358
rect 17316 18294 17368 18300
rect 16948 18284 17000 18290
rect 16948 18226 17000 18232
rect 16396 18216 16448 18222
rect 16396 18158 16448 18164
rect 16672 18216 16724 18222
rect 16672 18158 16724 18164
rect 16304 17536 16356 17542
rect 16304 17478 16356 17484
rect 16316 16522 16344 17478
rect 16304 16516 16356 16522
rect 16304 16458 16356 16464
rect 16408 16454 16436 18158
rect 16486 17640 16542 17649
rect 16486 17575 16488 17584
rect 16540 17575 16542 17584
rect 16488 17546 16540 17552
rect 16396 16448 16448 16454
rect 16396 16390 16448 16396
rect 16212 15156 16264 15162
rect 16212 15098 16264 15104
rect 16210 15056 16266 15065
rect 16210 14991 16212 15000
rect 16264 14991 16266 15000
rect 16212 14962 16264 14968
rect 16408 14958 16436 16390
rect 16684 16182 16712 18158
rect 17052 16946 17080 18294
rect 17592 17876 17644 17882
rect 17592 17818 17644 17824
rect 17604 17202 17632 17818
rect 17592 17196 17644 17202
rect 17592 17138 17644 17144
rect 17224 17128 17276 17134
rect 17224 17070 17276 17076
rect 16960 16918 17080 16946
rect 16856 16788 16908 16794
rect 16856 16730 16908 16736
rect 16764 16516 16816 16522
rect 16764 16458 16816 16464
rect 16672 16176 16724 16182
rect 16672 16118 16724 16124
rect 16488 16108 16540 16114
rect 16488 16050 16540 16056
rect 16500 15026 16528 16050
rect 16776 15162 16804 16458
rect 16868 16046 16896 16730
rect 16960 16250 16988 16918
rect 17236 16794 17264 17070
rect 17500 16992 17552 16998
rect 17500 16934 17552 16940
rect 17224 16788 17276 16794
rect 17224 16730 17276 16736
rect 17236 16590 17264 16730
rect 17316 16652 17368 16658
rect 17316 16594 17368 16600
rect 17224 16584 17276 16590
rect 17224 16526 17276 16532
rect 16948 16244 17000 16250
rect 16948 16186 17000 16192
rect 16856 16040 16908 16046
rect 16856 15982 16908 15988
rect 16764 15156 16816 15162
rect 16764 15098 16816 15104
rect 16488 15020 16540 15026
rect 16488 14962 16540 14968
rect 16396 14952 16448 14958
rect 16396 14894 16448 14900
rect 16500 14550 16528 14962
rect 16776 14618 16804 15098
rect 16960 15065 16988 16186
rect 17328 16182 17356 16594
rect 17316 16176 17368 16182
rect 17316 16118 17368 16124
rect 17130 15464 17186 15473
rect 17130 15399 17186 15408
rect 17144 15366 17172 15399
rect 17132 15360 17184 15366
rect 17132 15302 17184 15308
rect 16946 15056 17002 15065
rect 16856 15020 16908 15026
rect 16946 14991 17002 15000
rect 16856 14962 16908 14968
rect 16764 14612 16816 14618
rect 16764 14554 16816 14560
rect 16396 14544 16448 14550
rect 16396 14486 16448 14492
rect 16488 14544 16540 14550
rect 16488 14486 16540 14492
rect 16028 14476 16080 14482
rect 16028 14418 16080 14424
rect 16120 14476 16172 14482
rect 16120 14418 16172 14424
rect 15936 14340 15988 14346
rect 15936 14282 15988 14288
rect 15844 14000 15896 14006
rect 15844 13942 15896 13948
rect 15948 13682 15976 14282
rect 16040 13802 16068 14418
rect 16028 13796 16080 13802
rect 16028 13738 16080 13744
rect 15948 13654 16068 13682
rect 16040 13394 16068 13654
rect 16132 13394 16160 14418
rect 16408 14346 16436 14486
rect 16396 14340 16448 14346
rect 16396 14282 16448 14288
rect 16500 13818 16528 14486
rect 16672 13864 16724 13870
rect 16396 13796 16448 13802
rect 16500 13790 16620 13818
rect 16672 13806 16724 13812
rect 16396 13738 16448 13744
rect 16028 13388 16080 13394
rect 16028 13330 16080 13336
rect 16120 13388 16172 13394
rect 16120 13330 16172 13336
rect 15620 13280 15700 13308
rect 15752 13320 15804 13326
rect 15568 13262 15620 13268
rect 15752 13262 15804 13268
rect 15936 13184 15988 13190
rect 15936 13126 15988 13132
rect 15660 12980 15712 12986
rect 15660 12922 15712 12928
rect 15568 12776 15620 12782
rect 15568 12718 15620 12724
rect 15580 12238 15608 12718
rect 15568 12232 15620 12238
rect 15568 12174 15620 12180
rect 15672 11354 15700 12922
rect 15948 12918 15976 13126
rect 15936 12912 15988 12918
rect 15936 12854 15988 12860
rect 15844 12844 15896 12850
rect 15844 12786 15896 12792
rect 15856 11898 15884 12786
rect 15844 11892 15896 11898
rect 15844 11834 15896 11840
rect 15476 11348 15528 11354
rect 15476 11290 15528 11296
rect 15660 11348 15712 11354
rect 15660 11290 15712 11296
rect 15292 10668 15344 10674
rect 15292 10610 15344 10616
rect 15200 10464 15252 10470
rect 15200 10406 15252 10412
rect 14846 10364 15154 10384
rect 14846 10362 14852 10364
rect 14908 10362 14932 10364
rect 14988 10362 15012 10364
rect 15068 10362 15092 10364
rect 15148 10362 15154 10364
rect 14908 10310 14910 10362
rect 15090 10310 15092 10362
rect 14846 10308 14852 10310
rect 14908 10308 14932 10310
rect 14988 10308 15012 10310
rect 15068 10308 15092 10310
rect 15148 10308 15154 10310
rect 14846 10288 15154 10308
rect 15488 10062 15516 11290
rect 15660 11212 15712 11218
rect 15660 11154 15712 11160
rect 14740 10056 14792 10062
rect 14740 9998 14792 10004
rect 15476 10056 15528 10062
rect 15476 9998 15528 10004
rect 14648 9988 14700 9994
rect 14648 9930 14700 9936
rect 14752 9722 14780 9998
rect 15488 9926 15516 9998
rect 15384 9920 15436 9926
rect 15384 9862 15436 9868
rect 15476 9920 15528 9926
rect 15476 9862 15528 9868
rect 14740 9716 14792 9722
rect 14740 9658 14792 9664
rect 14846 9276 15154 9296
rect 14846 9274 14852 9276
rect 14908 9274 14932 9276
rect 14988 9274 15012 9276
rect 15068 9274 15092 9276
rect 15148 9274 15154 9276
rect 14908 9222 14910 9274
rect 15090 9222 15092 9274
rect 14846 9220 14852 9222
rect 14908 9220 14932 9222
rect 14988 9220 15012 9222
rect 15068 9220 15092 9222
rect 15148 9220 15154 9222
rect 14846 9200 15154 9220
rect 15292 9104 15344 9110
rect 15292 9046 15344 9052
rect 15200 9036 15252 9042
rect 15200 8978 15252 8984
rect 15212 8906 15240 8978
rect 15200 8900 15252 8906
rect 15200 8842 15252 8848
rect 15200 8492 15252 8498
rect 15200 8434 15252 8440
rect 14740 8424 14792 8430
rect 14740 8366 14792 8372
rect 14648 7336 14700 7342
rect 14648 7278 14700 7284
rect 14660 6390 14688 7278
rect 14752 6798 14780 8366
rect 14846 8188 15154 8208
rect 14846 8186 14852 8188
rect 14908 8186 14932 8188
rect 14988 8186 15012 8188
rect 15068 8186 15092 8188
rect 15148 8186 15154 8188
rect 14908 8134 14910 8186
rect 15090 8134 15092 8186
rect 14846 8132 14852 8134
rect 14908 8132 14932 8134
rect 14988 8132 15012 8134
rect 15068 8132 15092 8134
rect 15148 8132 15154 8134
rect 14846 8112 15154 8132
rect 15212 8090 15240 8434
rect 15304 8090 15332 9046
rect 15200 8084 15252 8090
rect 15200 8026 15252 8032
rect 15292 8084 15344 8090
rect 15292 8026 15344 8032
rect 14846 7100 15154 7120
rect 14846 7098 14852 7100
rect 14908 7098 14932 7100
rect 14988 7098 15012 7100
rect 15068 7098 15092 7100
rect 15148 7098 15154 7100
rect 14908 7046 14910 7098
rect 15090 7046 15092 7098
rect 14846 7044 14852 7046
rect 14908 7044 14932 7046
rect 14988 7044 15012 7046
rect 15068 7044 15092 7046
rect 15148 7044 15154 7046
rect 14846 7024 15154 7044
rect 14740 6792 14792 6798
rect 14740 6734 14792 6740
rect 14648 6384 14700 6390
rect 14648 6326 14700 6332
rect 14846 6012 15154 6032
rect 14846 6010 14852 6012
rect 14908 6010 14932 6012
rect 14988 6010 15012 6012
rect 15068 6010 15092 6012
rect 15148 6010 15154 6012
rect 14908 5958 14910 6010
rect 15090 5958 15092 6010
rect 14846 5956 14852 5958
rect 14908 5956 14932 5958
rect 14988 5956 15012 5958
rect 15068 5956 15092 5958
rect 15148 5956 15154 5958
rect 14846 5936 15154 5956
rect 15396 5846 15424 9862
rect 15568 8288 15620 8294
rect 15568 8230 15620 8236
rect 15580 7954 15608 8230
rect 15568 7948 15620 7954
rect 15568 7890 15620 7896
rect 15476 7472 15528 7478
rect 15476 7414 15528 7420
rect 15488 7002 15516 7414
rect 15476 6996 15528 7002
rect 15476 6938 15528 6944
rect 15488 6322 15516 6938
rect 15476 6316 15528 6322
rect 15476 6258 15528 6264
rect 15384 5840 15436 5846
rect 15384 5782 15436 5788
rect 14556 5636 14608 5642
rect 14556 5578 14608 5584
rect 14280 5568 14332 5574
rect 14280 5510 14332 5516
rect 14292 5234 14320 5510
rect 14004 5228 14056 5234
rect 14004 5170 14056 5176
rect 14280 5228 14332 5234
rect 14280 5170 14332 5176
rect 13912 5160 13964 5166
rect 13912 5102 13964 5108
rect 13452 5024 13504 5030
rect 13452 4966 13504 4972
rect 13544 5024 13596 5030
rect 13544 4966 13596 4972
rect 13360 4752 13412 4758
rect 13360 4694 13412 4700
rect 13176 4616 13228 4622
rect 13176 4558 13228 4564
rect 13188 4298 13216 4558
rect 13188 4270 13308 4298
rect 13176 4140 13228 4146
rect 13176 4082 13228 4088
rect 13084 3732 13136 3738
rect 13084 3674 13136 3680
rect 13188 3602 13216 4082
rect 13280 3942 13308 4270
rect 13268 3936 13320 3942
rect 13268 3878 13320 3884
rect 13280 3670 13308 3878
rect 13268 3664 13320 3670
rect 13268 3606 13320 3612
rect 13176 3596 13228 3602
rect 13176 3538 13228 3544
rect 12624 3528 12676 3534
rect 12624 3470 12676 3476
rect 13188 3194 13216 3538
rect 11980 3188 12032 3194
rect 11980 3130 12032 3136
rect 13176 3188 13228 3194
rect 13176 3130 13228 3136
rect 10968 2984 11020 2990
rect 10968 2926 11020 2932
rect 13280 2922 13308 3606
rect 13464 3534 13492 4966
rect 13556 3602 13584 4966
rect 13728 3664 13780 3670
rect 13728 3606 13780 3612
rect 13544 3596 13596 3602
rect 13544 3538 13596 3544
rect 13452 3528 13504 3534
rect 13452 3470 13504 3476
rect 13740 3058 13768 3606
rect 14016 3466 14044 5170
rect 14568 5166 14596 5578
rect 15292 5296 15344 5302
rect 15292 5238 15344 5244
rect 14556 5160 14608 5166
rect 14556 5102 14608 5108
rect 14188 5024 14240 5030
rect 14188 4966 14240 4972
rect 14096 4616 14148 4622
rect 14096 4558 14148 4564
rect 14108 4282 14136 4558
rect 14096 4276 14148 4282
rect 14096 4218 14148 4224
rect 14200 4214 14228 4966
rect 14568 4622 14596 5102
rect 14740 5024 14792 5030
rect 14740 4966 14792 4972
rect 14752 4690 14780 4966
rect 14846 4924 15154 4944
rect 14846 4922 14852 4924
rect 14908 4922 14932 4924
rect 14988 4922 15012 4924
rect 15068 4922 15092 4924
rect 15148 4922 15154 4924
rect 14908 4870 14910 4922
rect 15090 4870 15092 4922
rect 14846 4868 14852 4870
rect 14908 4868 14932 4870
rect 14988 4868 15012 4870
rect 15068 4868 15092 4870
rect 15148 4868 15154 4870
rect 14846 4848 15154 4868
rect 14740 4684 14792 4690
rect 14740 4626 14792 4632
rect 14556 4616 14608 4622
rect 14556 4558 14608 4564
rect 15304 4554 15332 5238
rect 15396 5030 15424 5782
rect 15384 5024 15436 5030
rect 15384 4966 15436 4972
rect 15292 4548 15344 4554
rect 15292 4490 15344 4496
rect 14188 4208 14240 4214
rect 14188 4150 14240 4156
rect 15384 4072 15436 4078
rect 15384 4014 15436 4020
rect 14846 3836 15154 3856
rect 14846 3834 14852 3836
rect 14908 3834 14932 3836
rect 14988 3834 15012 3836
rect 15068 3834 15092 3836
rect 15148 3834 15154 3836
rect 14908 3782 14910 3834
rect 15090 3782 15092 3834
rect 14846 3780 14852 3782
rect 14908 3780 14932 3782
rect 14988 3780 15012 3782
rect 15068 3780 15092 3782
rect 15148 3780 15154 3782
rect 14846 3760 15154 3780
rect 14004 3460 14056 3466
rect 14004 3402 14056 3408
rect 15396 3126 15424 4014
rect 15384 3120 15436 3126
rect 15384 3062 15436 3068
rect 13728 3052 13780 3058
rect 13728 2994 13780 3000
rect 13268 2916 13320 2922
rect 13268 2858 13320 2864
rect 1676 2848 1728 2854
rect 1676 2790 1728 2796
rect 5908 2848 5960 2854
rect 5908 2790 5960 2796
rect 1688 2378 1716 2790
rect 5582 2748 5890 2768
rect 5582 2746 5588 2748
rect 5644 2746 5668 2748
rect 5724 2746 5748 2748
rect 5804 2746 5828 2748
rect 5884 2746 5890 2748
rect 5644 2694 5646 2746
rect 5826 2694 5828 2746
rect 5582 2692 5588 2694
rect 5644 2692 5668 2694
rect 5724 2692 5748 2694
rect 5804 2692 5828 2694
rect 5884 2692 5890 2694
rect 5582 2672 5890 2692
rect 5920 2514 5948 2790
rect 14846 2748 15154 2768
rect 14846 2746 14852 2748
rect 14908 2746 14932 2748
rect 14988 2746 15012 2748
rect 15068 2746 15092 2748
rect 15148 2746 15154 2748
rect 14908 2694 14910 2746
rect 15090 2694 15092 2746
rect 14846 2692 14852 2694
rect 14908 2692 14932 2694
rect 14988 2692 15012 2694
rect 15068 2692 15092 2694
rect 15148 2692 15154 2694
rect 14846 2672 15154 2692
rect 5908 2508 5960 2514
rect 5908 2450 5960 2456
rect 3240 2440 3292 2446
rect 3240 2382 3292 2388
rect 6460 2440 6512 2446
rect 6460 2382 6512 2388
rect 12256 2440 12308 2446
rect 12256 2382 12308 2388
rect 1676 2372 1728 2378
rect 1676 2314 1728 2320
rect 18 0 74 800
rect 662 0 718 800
rect 1688 785 1716 2314
rect 2228 2304 2280 2310
rect 2228 2246 2280 2252
rect 2240 2145 2268 2246
rect 2226 2136 2282 2145
rect 2226 2071 2282 2080
rect 3252 800 3280 2382
rect 5172 2304 5224 2310
rect 5172 2246 5224 2252
rect 5184 800 5212 2246
rect 6472 800 6500 2382
rect 10214 2204 10522 2224
rect 10214 2202 10220 2204
rect 10276 2202 10300 2204
rect 10356 2202 10380 2204
rect 10436 2202 10460 2204
rect 10516 2202 10522 2204
rect 10276 2150 10278 2202
rect 10458 2150 10460 2202
rect 10214 2148 10220 2150
rect 10276 2148 10300 2150
rect 10356 2148 10380 2150
rect 10436 2148 10460 2150
rect 10516 2148 10522 2150
rect 10214 2128 10522 2148
rect 12268 800 12296 2382
rect 15672 2378 15700 11154
rect 15844 10464 15896 10470
rect 15844 10406 15896 10412
rect 15856 10130 15884 10406
rect 15844 10124 15896 10130
rect 15844 10066 15896 10072
rect 15856 9586 15884 10066
rect 15844 9580 15896 9586
rect 15844 9522 15896 9528
rect 15844 8628 15896 8634
rect 15844 8570 15896 8576
rect 15856 7410 15884 8570
rect 16040 7426 16068 13330
rect 16408 13326 16436 13738
rect 16592 13326 16620 13790
rect 16684 13462 16712 13806
rect 16776 13530 16804 14554
rect 16764 13524 16816 13530
rect 16764 13466 16816 13472
rect 16672 13456 16724 13462
rect 16672 13398 16724 13404
rect 16396 13320 16448 13326
rect 16396 13262 16448 13268
rect 16580 13320 16632 13326
rect 16580 13262 16632 13268
rect 16396 12912 16448 12918
rect 16396 12854 16448 12860
rect 16120 12640 16172 12646
rect 16120 12582 16172 12588
rect 16132 12238 16160 12582
rect 16408 12238 16436 12854
rect 16684 12850 16712 13398
rect 16868 13394 16896 14962
rect 16948 14408 17000 14414
rect 17040 14408 17092 14414
rect 16948 14350 17000 14356
rect 17038 14376 17040 14385
rect 17092 14376 17094 14385
rect 16856 13388 16908 13394
rect 16856 13330 16908 13336
rect 16960 12986 16988 14350
rect 17038 14311 17094 14320
rect 17040 13932 17092 13938
rect 17040 13874 17092 13880
rect 17052 13258 17080 13874
rect 17408 13320 17460 13326
rect 17408 13262 17460 13268
rect 17040 13252 17092 13258
rect 17040 13194 17092 13200
rect 17224 13184 17276 13190
rect 17224 13126 17276 13132
rect 16948 12980 17000 12986
rect 16948 12922 17000 12928
rect 16672 12844 16724 12850
rect 16672 12786 16724 12792
rect 16856 12776 16908 12782
rect 16856 12718 16908 12724
rect 16672 12708 16724 12714
rect 16672 12650 16724 12656
rect 16580 12640 16632 12646
rect 16580 12582 16632 12588
rect 16592 12442 16620 12582
rect 16580 12436 16632 12442
rect 16580 12378 16632 12384
rect 16120 12232 16172 12238
rect 16120 12174 16172 12180
rect 16396 12232 16448 12238
rect 16396 12174 16448 12180
rect 16580 12096 16632 12102
rect 16580 12038 16632 12044
rect 16592 11830 16620 12038
rect 16580 11824 16632 11830
rect 16580 11766 16632 11772
rect 16120 11552 16172 11558
rect 16120 11494 16172 11500
rect 16132 11082 16160 11494
rect 16304 11280 16356 11286
rect 16304 11222 16356 11228
rect 16120 11076 16172 11082
rect 16120 11018 16172 11024
rect 16132 8945 16160 11018
rect 16316 10198 16344 11222
rect 16684 10810 16712 12650
rect 16868 11286 16896 12718
rect 17236 12646 17264 13126
rect 17420 12986 17448 13262
rect 17408 12980 17460 12986
rect 17408 12922 17460 12928
rect 17512 12850 17540 16934
rect 17604 13433 17632 17138
rect 17788 16454 17816 18770
rect 17960 18760 18012 18766
rect 17960 18702 18012 18708
rect 18144 18760 18196 18766
rect 18144 18702 18196 18708
rect 17972 17202 18000 18702
rect 18052 18624 18104 18630
rect 18052 18566 18104 18572
rect 18064 18086 18092 18566
rect 18052 18080 18104 18086
rect 18052 18022 18104 18028
rect 17960 17196 18012 17202
rect 17960 17138 18012 17144
rect 18064 16454 18092 18022
rect 18156 17882 18184 18702
rect 18144 17876 18196 17882
rect 18144 17818 18196 17824
rect 18248 17542 18276 19722
rect 18800 19514 18828 20402
rect 19168 20058 19196 20402
rect 19260 20058 19288 20742
rect 19352 20602 19380 20946
rect 19904 20874 19932 21898
rect 19996 21554 20024 23054
rect 20272 22234 20300 23054
rect 20260 22228 20312 22234
rect 20260 22170 20312 22176
rect 20548 22030 20576 23258
rect 20916 22710 20944 23734
rect 21180 23520 21232 23526
rect 21180 23462 21232 23468
rect 20904 22704 20956 22710
rect 20904 22646 20956 22652
rect 20628 22636 20680 22642
rect 20628 22578 20680 22584
rect 20536 22024 20588 22030
rect 20536 21966 20588 21972
rect 20548 21690 20576 21966
rect 20536 21684 20588 21690
rect 20536 21626 20588 21632
rect 19984 21548 20036 21554
rect 19984 21490 20036 21496
rect 20168 21548 20220 21554
rect 20168 21490 20220 21496
rect 20260 21548 20312 21554
rect 20260 21490 20312 21496
rect 19984 21412 20036 21418
rect 19984 21354 20036 21360
rect 19892 20868 19944 20874
rect 19892 20810 19944 20816
rect 19478 20700 19786 20720
rect 19478 20698 19484 20700
rect 19540 20698 19564 20700
rect 19620 20698 19644 20700
rect 19700 20698 19724 20700
rect 19780 20698 19786 20700
rect 19540 20646 19542 20698
rect 19722 20646 19724 20698
rect 19478 20644 19484 20646
rect 19540 20644 19564 20646
rect 19620 20644 19644 20646
rect 19700 20644 19724 20646
rect 19780 20644 19786 20646
rect 19478 20624 19786 20644
rect 19340 20596 19392 20602
rect 19340 20538 19392 20544
rect 19996 20466 20024 21354
rect 20180 20602 20208 21490
rect 20272 21146 20300 21490
rect 20260 21140 20312 21146
rect 20260 21082 20312 21088
rect 20536 20868 20588 20874
rect 20536 20810 20588 20816
rect 20260 20800 20312 20806
rect 20260 20742 20312 20748
rect 20444 20800 20496 20806
rect 20444 20742 20496 20748
rect 20168 20596 20220 20602
rect 20168 20538 20220 20544
rect 19984 20460 20036 20466
rect 19984 20402 20036 20408
rect 20168 20460 20220 20466
rect 20168 20402 20220 20408
rect 19156 20052 19208 20058
rect 19156 19994 19208 20000
rect 19248 20052 19300 20058
rect 19248 19994 19300 20000
rect 19892 19916 19944 19922
rect 19892 19858 19944 19864
rect 19478 19612 19786 19632
rect 19478 19610 19484 19612
rect 19540 19610 19564 19612
rect 19620 19610 19644 19612
rect 19700 19610 19724 19612
rect 19780 19610 19786 19612
rect 19540 19558 19542 19610
rect 19722 19558 19724 19610
rect 19478 19556 19484 19558
rect 19540 19556 19564 19558
rect 19620 19556 19644 19558
rect 19700 19556 19724 19558
rect 19780 19556 19786 19558
rect 19478 19536 19786 19556
rect 18788 19508 18840 19514
rect 18788 19450 18840 19456
rect 19340 19440 19392 19446
rect 19340 19382 19392 19388
rect 19616 19440 19668 19446
rect 19616 19382 19668 19388
rect 19352 18970 19380 19382
rect 19628 19174 19656 19382
rect 19616 19168 19668 19174
rect 19616 19110 19668 19116
rect 19340 18964 19392 18970
rect 19340 18906 19392 18912
rect 19248 18692 19300 18698
rect 19248 18634 19300 18640
rect 18328 18624 18380 18630
rect 18328 18566 18380 18572
rect 18340 18290 18368 18566
rect 19260 18290 19288 18634
rect 19352 18358 19380 18906
rect 19628 18698 19656 19110
rect 19616 18692 19668 18698
rect 19616 18634 19668 18640
rect 19478 18524 19786 18544
rect 19478 18522 19484 18524
rect 19540 18522 19564 18524
rect 19620 18522 19644 18524
rect 19700 18522 19724 18524
rect 19780 18522 19786 18524
rect 19540 18470 19542 18522
rect 19722 18470 19724 18522
rect 19478 18468 19484 18470
rect 19540 18468 19564 18470
rect 19620 18468 19644 18470
rect 19700 18468 19724 18470
rect 19780 18468 19786 18470
rect 19478 18448 19786 18468
rect 19904 18426 19932 19858
rect 19892 18420 19944 18426
rect 19892 18362 19944 18368
rect 19340 18352 19392 18358
rect 19340 18294 19392 18300
rect 18328 18284 18380 18290
rect 18328 18226 18380 18232
rect 19248 18284 19300 18290
rect 19248 18226 19300 18232
rect 18604 17876 18656 17882
rect 18604 17818 18656 17824
rect 18616 17610 18644 17818
rect 19352 17746 19380 18294
rect 19340 17740 19392 17746
rect 19340 17682 19392 17688
rect 18512 17604 18564 17610
rect 18512 17546 18564 17552
rect 18604 17604 18656 17610
rect 18604 17546 18656 17552
rect 18236 17536 18288 17542
rect 18236 17478 18288 17484
rect 18248 17338 18276 17478
rect 18524 17338 18552 17546
rect 18236 17332 18288 17338
rect 18236 17274 18288 17280
rect 18512 17332 18564 17338
rect 18512 17274 18564 17280
rect 18326 17232 18382 17241
rect 18326 17167 18382 17176
rect 18340 16794 18368 17167
rect 18328 16788 18380 16794
rect 18328 16730 18380 16736
rect 17776 16448 17828 16454
rect 17776 16390 17828 16396
rect 18052 16448 18104 16454
rect 18052 16390 18104 16396
rect 18236 16448 18288 16454
rect 18236 16390 18288 16396
rect 17776 16244 17828 16250
rect 17776 16186 17828 16192
rect 17788 15910 17816 16186
rect 17868 16108 17920 16114
rect 17868 16050 17920 16056
rect 17776 15904 17828 15910
rect 17776 15846 17828 15852
rect 17788 15162 17816 15846
rect 17880 15570 17908 16050
rect 17868 15564 17920 15570
rect 17868 15506 17920 15512
rect 17776 15156 17828 15162
rect 17776 15098 17828 15104
rect 17682 15056 17738 15065
rect 17682 14991 17738 15000
rect 17866 15056 17922 15065
rect 17866 14991 17922 15000
rect 17696 14822 17724 14991
rect 17684 14816 17736 14822
rect 17684 14758 17736 14764
rect 17776 14544 17828 14550
rect 17776 14486 17828 14492
rect 17788 13938 17816 14486
rect 17880 14414 17908 14991
rect 18052 14816 18104 14822
rect 18052 14758 18104 14764
rect 18064 14618 18092 14758
rect 18052 14612 18104 14618
rect 18052 14554 18104 14560
rect 18064 14414 18092 14554
rect 17868 14408 17920 14414
rect 17868 14350 17920 14356
rect 18052 14408 18104 14414
rect 18052 14350 18104 14356
rect 17776 13932 17828 13938
rect 17776 13874 17828 13880
rect 17590 13424 17646 13433
rect 17590 13359 17646 13368
rect 17604 13326 17632 13359
rect 17592 13320 17644 13326
rect 17592 13262 17644 13268
rect 17500 12844 17552 12850
rect 17500 12786 17552 12792
rect 17224 12640 17276 12646
rect 17224 12582 17276 12588
rect 17316 12640 17368 12646
rect 17316 12582 17368 12588
rect 17236 12306 17264 12582
rect 17040 12300 17092 12306
rect 17040 12242 17092 12248
rect 17224 12300 17276 12306
rect 17224 12242 17276 12248
rect 17052 11762 17080 12242
rect 17328 12238 17356 12582
rect 17592 12368 17644 12374
rect 17592 12310 17644 12316
rect 17316 12232 17368 12238
rect 17316 12174 17368 12180
rect 17500 12232 17552 12238
rect 17500 12174 17552 12180
rect 17512 12073 17540 12174
rect 17498 12064 17554 12073
rect 17498 11999 17554 12008
rect 17040 11756 17092 11762
rect 17040 11698 17092 11704
rect 17052 11354 17080 11698
rect 17512 11354 17540 11999
rect 17040 11348 17092 11354
rect 17040 11290 17092 11296
rect 17500 11348 17552 11354
rect 17500 11290 17552 11296
rect 16856 11280 16908 11286
rect 16856 11222 16908 11228
rect 16672 10804 16724 10810
rect 16672 10746 16724 10752
rect 16304 10192 16356 10198
rect 16304 10134 16356 10140
rect 16316 9586 16344 10134
rect 16764 10056 16816 10062
rect 17512 10010 17540 11290
rect 16764 9998 16816 10004
rect 16580 9920 16632 9926
rect 16580 9862 16632 9868
rect 16304 9580 16356 9586
rect 16304 9522 16356 9528
rect 16316 9450 16344 9522
rect 16304 9444 16356 9450
rect 16304 9386 16356 9392
rect 16118 8936 16174 8945
rect 16118 8871 16174 8880
rect 16212 8560 16264 8566
rect 16212 8502 16264 8508
rect 16224 8090 16252 8502
rect 16212 8084 16264 8090
rect 16212 8026 16264 8032
rect 16488 8084 16540 8090
rect 16488 8026 16540 8032
rect 16500 7750 16528 8026
rect 16488 7744 16540 7750
rect 16488 7686 16540 7692
rect 16500 7478 16528 7686
rect 16488 7472 16540 7478
rect 15844 7404 15896 7410
rect 15844 7346 15896 7352
rect 15936 7404 15988 7410
rect 16040 7398 16160 7426
rect 16488 7414 16540 7420
rect 15936 7346 15988 7352
rect 15948 6458 15976 7346
rect 16028 7200 16080 7206
rect 16028 7142 16080 7148
rect 16040 6798 16068 7142
rect 16028 6792 16080 6798
rect 16028 6734 16080 6740
rect 15936 6452 15988 6458
rect 15936 6394 15988 6400
rect 16132 5370 16160 7398
rect 16592 5710 16620 9862
rect 16776 9722 16804 9998
rect 17236 9982 17540 10010
rect 17604 9994 17632 12310
rect 17776 12096 17828 12102
rect 17776 12038 17828 12044
rect 17788 11082 17816 12038
rect 17880 11898 17908 14350
rect 17960 13728 18012 13734
rect 17960 13670 18012 13676
rect 18144 13728 18196 13734
rect 18144 13670 18196 13676
rect 17972 13530 18000 13670
rect 17960 13524 18012 13530
rect 17960 13466 18012 13472
rect 17972 13258 18000 13466
rect 18052 13388 18104 13394
rect 18052 13330 18104 13336
rect 17960 13252 18012 13258
rect 17960 13194 18012 13200
rect 18064 12170 18092 13330
rect 18052 12164 18104 12170
rect 18052 12106 18104 12112
rect 17868 11892 17920 11898
rect 17868 11834 17920 11840
rect 18052 11688 18104 11694
rect 18052 11630 18104 11636
rect 18064 11150 18092 11630
rect 18052 11144 18104 11150
rect 18052 11086 18104 11092
rect 17776 11076 17828 11082
rect 17776 11018 17828 11024
rect 17684 10192 17736 10198
rect 17684 10134 17736 10140
rect 17592 9988 17644 9994
rect 16764 9716 16816 9722
rect 16764 9658 16816 9664
rect 16672 8900 16724 8906
rect 17040 8900 17092 8906
rect 16724 8860 17040 8888
rect 16672 8842 16724 8848
rect 17040 8842 17092 8848
rect 17052 8566 17080 8842
rect 17040 8560 17092 8566
rect 17040 8502 17092 8508
rect 16948 8356 17000 8362
rect 16948 8298 17000 8304
rect 16960 8090 16988 8298
rect 16948 8084 17000 8090
rect 16948 8026 17000 8032
rect 17040 7880 17092 7886
rect 17092 7840 17172 7868
rect 17040 7822 17092 7828
rect 17040 7404 17092 7410
rect 17040 7346 17092 7352
rect 16948 5840 17000 5846
rect 16948 5782 17000 5788
rect 16580 5704 16632 5710
rect 16578 5672 16580 5681
rect 16632 5672 16634 5681
rect 16578 5607 16634 5616
rect 16120 5364 16172 5370
rect 16120 5306 16172 5312
rect 16764 5296 16816 5302
rect 16764 5238 16816 5244
rect 16120 5024 16172 5030
rect 16120 4966 16172 4972
rect 16132 4622 16160 4966
rect 16120 4616 16172 4622
rect 16120 4558 16172 4564
rect 16672 4480 16724 4486
rect 16672 4422 16724 4428
rect 16684 4146 16712 4422
rect 16672 4140 16724 4146
rect 16672 4082 16724 4088
rect 16776 3534 16804 5238
rect 16960 5234 16988 5782
rect 16948 5228 17000 5234
rect 16948 5170 17000 5176
rect 17052 4214 17080 7346
rect 17144 6662 17172 7840
rect 17132 6656 17184 6662
rect 17132 6598 17184 6604
rect 17144 6254 17172 6598
rect 17132 6248 17184 6254
rect 17132 6190 17184 6196
rect 17236 6100 17264 9982
rect 17592 9930 17644 9936
rect 17604 9586 17632 9930
rect 17696 9654 17724 10134
rect 17960 9920 18012 9926
rect 17960 9862 18012 9868
rect 17684 9648 17736 9654
rect 17684 9590 17736 9596
rect 17316 9580 17368 9586
rect 17316 9522 17368 9528
rect 17408 9580 17460 9586
rect 17592 9580 17644 9586
rect 17408 9522 17460 9528
rect 17512 9540 17592 9568
rect 17328 9178 17356 9522
rect 17316 9172 17368 9178
rect 17316 9114 17368 9120
rect 17420 8634 17448 9522
rect 17408 8628 17460 8634
rect 17408 8570 17460 8576
rect 17316 7744 17368 7750
rect 17316 7686 17368 7692
rect 17328 6866 17356 7686
rect 17512 7546 17540 9540
rect 17592 9522 17644 9528
rect 17776 9376 17828 9382
rect 17776 9318 17828 9324
rect 17788 8974 17816 9318
rect 17592 8968 17644 8974
rect 17592 8910 17644 8916
rect 17776 8968 17828 8974
rect 17776 8910 17828 8916
rect 17604 8430 17632 8910
rect 17868 8832 17920 8838
rect 17868 8774 17920 8780
rect 17880 8566 17908 8774
rect 17868 8560 17920 8566
rect 17868 8502 17920 8508
rect 17592 8424 17644 8430
rect 17592 8366 17644 8372
rect 17408 7540 17460 7546
rect 17408 7482 17460 7488
rect 17500 7540 17552 7546
rect 17500 7482 17552 7488
rect 17420 7002 17448 7482
rect 17604 7410 17632 8366
rect 17880 7886 17908 8502
rect 17868 7880 17920 7886
rect 17868 7822 17920 7828
rect 17500 7404 17552 7410
rect 17500 7346 17552 7352
rect 17592 7404 17644 7410
rect 17592 7346 17644 7352
rect 17408 6996 17460 7002
rect 17408 6938 17460 6944
rect 17512 6934 17540 7346
rect 17500 6928 17552 6934
rect 17500 6870 17552 6876
rect 17316 6860 17368 6866
rect 17316 6802 17368 6808
rect 17500 6656 17552 6662
rect 17500 6598 17552 6604
rect 17512 6322 17540 6598
rect 17500 6316 17552 6322
rect 17500 6258 17552 6264
rect 17408 6180 17460 6186
rect 17408 6122 17460 6128
rect 17144 6072 17264 6100
rect 17040 4208 17092 4214
rect 17040 4150 17092 4156
rect 16948 3936 17000 3942
rect 16948 3878 17000 3884
rect 16764 3528 16816 3534
rect 16764 3470 16816 3476
rect 16960 3466 16988 3878
rect 16948 3460 17000 3466
rect 16948 3402 17000 3408
rect 17144 2774 17172 6072
rect 17420 5574 17448 6122
rect 17408 5568 17460 5574
rect 17408 5510 17460 5516
rect 17420 4826 17448 5510
rect 17604 5302 17632 7346
rect 17776 6792 17828 6798
rect 17776 6734 17828 6740
rect 17788 6254 17816 6734
rect 17972 6458 18000 9862
rect 18064 9586 18092 11086
rect 18156 9654 18184 13670
rect 18248 12209 18276 16390
rect 18340 16114 18368 16730
rect 18420 16516 18472 16522
rect 18420 16458 18472 16464
rect 18328 16108 18380 16114
rect 18328 16050 18380 16056
rect 18340 14958 18368 16050
rect 18432 15502 18460 16458
rect 18420 15496 18472 15502
rect 18420 15438 18472 15444
rect 18328 14952 18380 14958
rect 18328 14894 18380 14900
rect 18340 14482 18368 14894
rect 18512 14816 18564 14822
rect 18512 14758 18564 14764
rect 18328 14476 18380 14482
rect 18328 14418 18380 14424
rect 18340 14006 18368 14418
rect 18524 14414 18552 14758
rect 18616 14550 18644 17546
rect 19352 17202 19380 17682
rect 19904 17678 19932 18362
rect 19996 17898 20024 20402
rect 20076 19984 20128 19990
rect 20076 19926 20128 19932
rect 20088 19496 20116 19926
rect 20180 19718 20208 20402
rect 20272 19922 20300 20742
rect 20456 20534 20484 20742
rect 20444 20528 20496 20534
rect 20444 20470 20496 20476
rect 20548 20398 20576 20810
rect 20536 20392 20588 20398
rect 20536 20334 20588 20340
rect 20640 19938 20668 22578
rect 21192 22094 21220 23462
rect 21456 22976 21508 22982
rect 21456 22918 21508 22924
rect 21364 22636 21416 22642
rect 21364 22578 21416 22584
rect 21376 22234 21404 22578
rect 21364 22228 21416 22234
rect 21364 22170 21416 22176
rect 21100 22066 21220 22094
rect 20904 21344 20956 21350
rect 20904 21286 20956 21292
rect 20916 20466 20944 21286
rect 20904 20460 20956 20466
rect 20904 20402 20956 20408
rect 20260 19916 20312 19922
rect 20260 19858 20312 19864
rect 20364 19910 20668 19938
rect 20272 19786 20300 19858
rect 20260 19780 20312 19786
rect 20260 19722 20312 19728
rect 20168 19712 20220 19718
rect 20168 19654 20220 19660
rect 20088 19468 20300 19496
rect 20076 19372 20128 19378
rect 20076 19314 20128 19320
rect 20088 18630 20116 19314
rect 20272 18766 20300 19468
rect 20260 18760 20312 18766
rect 20260 18702 20312 18708
rect 20168 18692 20220 18698
rect 20168 18634 20220 18640
rect 20076 18624 20128 18630
rect 20076 18566 20128 18572
rect 20180 18426 20208 18634
rect 20168 18420 20220 18426
rect 20168 18362 20220 18368
rect 19996 17870 20208 17898
rect 19984 17740 20036 17746
rect 19984 17682 20036 17688
rect 19892 17672 19944 17678
rect 19892 17614 19944 17620
rect 19478 17436 19786 17456
rect 19478 17434 19484 17436
rect 19540 17434 19564 17436
rect 19620 17434 19644 17436
rect 19700 17434 19724 17436
rect 19780 17434 19786 17436
rect 19540 17382 19542 17434
rect 19722 17382 19724 17434
rect 19478 17380 19484 17382
rect 19540 17380 19564 17382
rect 19620 17380 19644 17382
rect 19700 17380 19724 17382
rect 19780 17380 19786 17382
rect 19478 17360 19786 17380
rect 18696 17196 18748 17202
rect 18696 17138 18748 17144
rect 19340 17196 19392 17202
rect 19340 17138 19392 17144
rect 18708 16454 18736 17138
rect 19616 17060 19668 17066
rect 19616 17002 19668 17008
rect 19064 16992 19116 16998
rect 19064 16934 19116 16940
rect 19524 16992 19576 16998
rect 19524 16934 19576 16940
rect 19076 16522 19104 16934
rect 19536 16794 19564 16934
rect 19628 16794 19656 17002
rect 19248 16788 19300 16794
rect 19248 16730 19300 16736
rect 19524 16788 19576 16794
rect 19524 16730 19576 16736
rect 19616 16788 19668 16794
rect 19616 16730 19668 16736
rect 19260 16590 19288 16730
rect 19248 16584 19300 16590
rect 19248 16526 19300 16532
rect 19064 16516 19116 16522
rect 19064 16458 19116 16464
rect 18696 16448 18748 16454
rect 18696 16390 18748 16396
rect 18604 14544 18656 14550
rect 18604 14486 18656 14492
rect 18512 14408 18564 14414
rect 18512 14350 18564 14356
rect 18420 14272 18472 14278
rect 18420 14214 18472 14220
rect 18328 14000 18380 14006
rect 18328 13942 18380 13948
rect 18432 13938 18460 14214
rect 18420 13932 18472 13938
rect 18420 13874 18472 13880
rect 18432 13326 18460 13874
rect 18420 13320 18472 13326
rect 18420 13262 18472 13268
rect 18328 13184 18380 13190
rect 18328 13126 18380 13132
rect 18234 12200 18290 12209
rect 18234 12135 18290 12144
rect 18144 9648 18196 9654
rect 18144 9590 18196 9596
rect 18052 9580 18104 9586
rect 18052 9522 18104 9528
rect 18248 9382 18276 12135
rect 18340 10742 18368 13126
rect 18524 11558 18552 14350
rect 18604 13728 18656 13734
rect 18604 13670 18656 13676
rect 18616 13326 18644 13670
rect 18604 13320 18656 13326
rect 18604 13262 18656 13268
rect 18512 11552 18564 11558
rect 18512 11494 18564 11500
rect 18328 10736 18380 10742
rect 18328 10678 18380 10684
rect 18328 10056 18380 10062
rect 18328 9998 18380 10004
rect 18236 9376 18288 9382
rect 18236 9318 18288 9324
rect 18248 8974 18276 9318
rect 18236 8968 18288 8974
rect 18236 8910 18288 8916
rect 18340 8090 18368 9998
rect 18708 9674 18736 16390
rect 18788 16108 18840 16114
rect 18788 16050 18840 16056
rect 18800 15858 18828 16050
rect 18800 15830 19012 15858
rect 18788 14884 18840 14890
rect 18788 14826 18840 14832
rect 18800 14550 18828 14826
rect 18984 14822 19012 15830
rect 19076 14890 19104 16458
rect 19892 16448 19944 16454
rect 19892 16390 19944 16396
rect 19478 16348 19786 16368
rect 19478 16346 19484 16348
rect 19540 16346 19564 16348
rect 19620 16346 19644 16348
rect 19700 16346 19724 16348
rect 19780 16346 19786 16348
rect 19540 16294 19542 16346
rect 19722 16294 19724 16346
rect 19478 16292 19484 16294
rect 19540 16292 19564 16294
rect 19620 16292 19644 16294
rect 19700 16292 19724 16294
rect 19780 16292 19786 16294
rect 19338 16280 19394 16289
rect 19156 16244 19208 16250
rect 19478 16272 19786 16292
rect 19338 16215 19340 16224
rect 19156 16186 19208 16192
rect 19392 16215 19394 16224
rect 19340 16186 19392 16192
rect 19168 16114 19196 16186
rect 19904 16114 19932 16390
rect 19156 16108 19208 16114
rect 19156 16050 19208 16056
rect 19892 16108 19944 16114
rect 19892 16050 19944 16056
rect 19432 15972 19484 15978
rect 19432 15914 19484 15920
rect 19444 15570 19472 15914
rect 19892 15904 19944 15910
rect 19892 15846 19944 15852
rect 19432 15564 19484 15570
rect 19352 15524 19432 15552
rect 19352 15026 19380 15524
rect 19432 15506 19484 15512
rect 19478 15260 19786 15280
rect 19478 15258 19484 15260
rect 19540 15258 19564 15260
rect 19620 15258 19644 15260
rect 19700 15258 19724 15260
rect 19780 15258 19786 15260
rect 19540 15206 19542 15258
rect 19722 15206 19724 15258
rect 19478 15204 19484 15206
rect 19540 15204 19564 15206
rect 19620 15204 19644 15206
rect 19700 15204 19724 15206
rect 19780 15204 19786 15206
rect 19478 15184 19786 15204
rect 19800 15088 19852 15094
rect 19798 15056 19800 15065
rect 19852 15056 19854 15065
rect 19340 15020 19392 15026
rect 19798 14991 19854 15000
rect 19340 14962 19392 14968
rect 19064 14884 19116 14890
rect 19064 14826 19116 14832
rect 18972 14816 19024 14822
rect 18972 14758 19024 14764
rect 18880 14612 18932 14618
rect 18880 14554 18932 14560
rect 18788 14544 18840 14550
rect 18788 14486 18840 14492
rect 18892 14278 18920 14554
rect 18880 14272 18932 14278
rect 18880 14214 18932 14220
rect 18892 14006 18920 14214
rect 18880 14000 18932 14006
rect 18880 13942 18932 13948
rect 18984 12986 19012 14758
rect 19076 14346 19104 14826
rect 19352 14482 19380 14962
rect 19524 14612 19576 14618
rect 19444 14572 19524 14600
rect 19340 14476 19392 14482
rect 19340 14418 19392 14424
rect 19248 14408 19300 14414
rect 19444 14362 19472 14572
rect 19904 14600 19932 15846
rect 19996 14618 20024 17682
rect 20180 16590 20208 17870
rect 20364 17746 20392 19910
rect 20628 19848 20680 19854
rect 20628 19790 20680 19796
rect 20536 19712 20588 19718
rect 20536 19654 20588 19660
rect 20444 19508 20496 19514
rect 20444 19450 20496 19456
rect 20456 18358 20484 19450
rect 20548 18630 20576 19654
rect 20640 19378 20668 19790
rect 21100 19718 21128 22066
rect 21468 22030 21496 22918
rect 21456 22024 21508 22030
rect 21456 21966 21508 21972
rect 21272 21344 21324 21350
rect 21272 21286 21324 21292
rect 21284 20942 21312 21286
rect 21272 20936 21324 20942
rect 21272 20878 21324 20884
rect 22100 19916 22152 19922
rect 22100 19858 22152 19864
rect 21732 19780 21784 19786
rect 21732 19722 21784 19728
rect 21088 19712 21140 19718
rect 21086 19680 21088 19689
rect 21140 19680 21142 19689
rect 21086 19615 21142 19624
rect 21744 19378 21772 19722
rect 20628 19372 20680 19378
rect 20628 19314 20680 19320
rect 20812 19372 20864 19378
rect 20812 19314 20864 19320
rect 21732 19372 21784 19378
rect 22112 19360 22140 19858
rect 22304 19372 22356 19378
rect 22112 19332 22304 19360
rect 21732 19314 21784 19320
rect 22304 19314 22356 19320
rect 20640 18970 20668 19314
rect 20720 19168 20772 19174
rect 20720 19110 20772 19116
rect 20732 18970 20760 19110
rect 20628 18964 20680 18970
rect 20628 18906 20680 18912
rect 20720 18964 20772 18970
rect 20720 18906 20772 18912
rect 20720 18760 20772 18766
rect 20720 18702 20772 18708
rect 20628 18692 20680 18698
rect 20628 18634 20680 18640
rect 20536 18624 20588 18630
rect 20536 18566 20588 18572
rect 20444 18352 20496 18358
rect 20444 18294 20496 18300
rect 20548 18154 20576 18566
rect 20640 18154 20668 18634
rect 20732 18358 20760 18702
rect 20720 18352 20772 18358
rect 20720 18294 20772 18300
rect 20824 18290 20852 19314
rect 20904 19304 20956 19310
rect 20904 19246 20956 19252
rect 20916 18358 20944 19246
rect 21456 19168 21508 19174
rect 21456 19110 21508 19116
rect 21468 18766 21496 19110
rect 22388 18970 22416 26930
rect 22848 23866 22876 27270
rect 23492 27130 23520 27270
rect 23480 27124 23532 27130
rect 23480 27066 23532 27072
rect 24032 26988 24084 26994
rect 24032 26930 24084 26936
rect 24044 26234 24072 26930
rect 24110 26684 24418 26704
rect 24110 26682 24116 26684
rect 24172 26682 24196 26684
rect 24252 26682 24276 26684
rect 24332 26682 24356 26684
rect 24412 26682 24418 26684
rect 24172 26630 24174 26682
rect 24354 26630 24356 26682
rect 24110 26628 24116 26630
rect 24172 26628 24196 26630
rect 24252 26628 24276 26630
rect 24332 26628 24356 26630
rect 24412 26628 24418 26630
rect 24110 26608 24418 26628
rect 23952 26206 24072 26234
rect 22836 23860 22888 23866
rect 22836 23802 22888 23808
rect 22468 20868 22520 20874
rect 22468 20810 22520 20816
rect 22376 18964 22428 18970
rect 22376 18906 22428 18912
rect 21824 18896 21876 18902
rect 21824 18838 21876 18844
rect 21180 18760 21232 18766
rect 21180 18702 21232 18708
rect 21456 18760 21508 18766
rect 21456 18702 21508 18708
rect 20904 18352 20956 18358
rect 20904 18294 20956 18300
rect 20812 18284 20864 18290
rect 20812 18226 20864 18232
rect 20536 18148 20588 18154
rect 20536 18090 20588 18096
rect 20628 18148 20680 18154
rect 20628 18090 20680 18096
rect 20444 18080 20496 18086
rect 20444 18022 20496 18028
rect 20352 17740 20404 17746
rect 20352 17682 20404 17688
rect 20260 17536 20312 17542
rect 20260 17478 20312 17484
rect 20272 17270 20300 17478
rect 20260 17264 20312 17270
rect 20260 17206 20312 17212
rect 20352 16992 20404 16998
rect 20456 16946 20484 18022
rect 20640 17814 20668 18090
rect 20720 18080 20772 18086
rect 20720 18022 20772 18028
rect 20732 17814 20760 18022
rect 20628 17808 20680 17814
rect 20628 17750 20680 17756
rect 20720 17808 20772 17814
rect 20720 17750 20772 17756
rect 20824 17490 20852 18226
rect 20916 17678 20944 18294
rect 21088 18284 21140 18290
rect 21088 18226 21140 18232
rect 20904 17672 20956 17678
rect 20904 17614 20956 17620
rect 20732 17462 20852 17490
rect 20732 16998 20760 17462
rect 21100 17338 21128 18226
rect 21088 17332 21140 17338
rect 21088 17274 21140 17280
rect 20404 16940 20484 16946
rect 20352 16934 20484 16940
rect 20720 16992 20772 16998
rect 20720 16934 20772 16940
rect 20364 16918 20484 16934
rect 20260 16652 20312 16658
rect 20260 16594 20312 16600
rect 20168 16584 20220 16590
rect 20168 16526 20220 16532
rect 20076 16108 20128 16114
rect 20076 16050 20128 16056
rect 20088 15502 20116 16050
rect 20076 15496 20128 15502
rect 20076 15438 20128 15444
rect 19576 14572 19932 14600
rect 19984 14612 20036 14618
rect 19524 14554 19576 14560
rect 19984 14554 20036 14560
rect 19248 14350 19300 14356
rect 19064 14340 19116 14346
rect 19064 14282 19116 14288
rect 19260 14074 19288 14350
rect 19352 14334 19472 14362
rect 19248 14068 19300 14074
rect 19248 14010 19300 14016
rect 19248 13320 19300 13326
rect 19248 13262 19300 13268
rect 19260 12986 19288 13262
rect 18972 12980 19024 12986
rect 18972 12922 19024 12928
rect 19248 12980 19300 12986
rect 19248 12922 19300 12928
rect 19352 12782 19380 14334
rect 19478 14172 19786 14192
rect 19478 14170 19484 14172
rect 19540 14170 19564 14172
rect 19620 14170 19644 14172
rect 19700 14170 19724 14172
rect 19780 14170 19786 14172
rect 19540 14118 19542 14170
rect 19722 14118 19724 14170
rect 19478 14116 19484 14118
rect 19540 14116 19564 14118
rect 19620 14116 19644 14118
rect 19700 14116 19724 14118
rect 19780 14116 19786 14118
rect 19478 14096 19786 14116
rect 19984 13932 20036 13938
rect 19984 13874 20036 13880
rect 19892 13320 19944 13326
rect 19892 13262 19944 13268
rect 19478 13084 19786 13104
rect 19478 13082 19484 13084
rect 19540 13082 19564 13084
rect 19620 13082 19644 13084
rect 19700 13082 19724 13084
rect 19780 13082 19786 13084
rect 19540 13030 19542 13082
rect 19722 13030 19724 13082
rect 19478 13028 19484 13030
rect 19540 13028 19564 13030
rect 19620 13028 19644 13030
rect 19700 13028 19724 13030
rect 19780 13028 19786 13030
rect 19478 13008 19786 13028
rect 18880 12776 18932 12782
rect 18880 12718 18932 12724
rect 19340 12776 19392 12782
rect 19340 12718 19392 12724
rect 18892 12646 18920 12718
rect 18880 12640 18932 12646
rect 18880 12582 18932 12588
rect 19340 12640 19392 12646
rect 19340 12582 19392 12588
rect 19352 12102 19380 12582
rect 19904 12170 19932 13262
rect 19996 12238 20024 13874
rect 20088 13530 20116 15438
rect 20180 14414 20208 16526
rect 20168 14408 20220 14414
rect 20168 14350 20220 14356
rect 20076 13524 20128 13530
rect 20076 13466 20128 13472
rect 20168 12844 20220 12850
rect 20168 12786 20220 12792
rect 20076 12776 20128 12782
rect 20076 12718 20128 12724
rect 19984 12232 20036 12238
rect 19984 12174 20036 12180
rect 19892 12164 19944 12170
rect 19892 12106 19944 12112
rect 19340 12096 19392 12102
rect 19340 12038 19392 12044
rect 18972 11552 19024 11558
rect 18972 11494 19024 11500
rect 19156 11552 19208 11558
rect 19156 11494 19208 11500
rect 18984 11082 19012 11494
rect 18972 11076 19024 11082
rect 18972 11018 19024 11024
rect 19168 10062 19196 11494
rect 19248 11144 19300 11150
rect 19248 11086 19300 11092
rect 19260 10810 19288 11086
rect 19248 10804 19300 10810
rect 19248 10746 19300 10752
rect 19260 10130 19288 10746
rect 19352 10554 19380 12038
rect 19478 11996 19786 12016
rect 19478 11994 19484 11996
rect 19540 11994 19564 11996
rect 19620 11994 19644 11996
rect 19700 11994 19724 11996
rect 19780 11994 19786 11996
rect 19540 11942 19542 11994
rect 19722 11942 19724 11994
rect 19478 11940 19484 11942
rect 19540 11940 19564 11942
rect 19620 11940 19644 11942
rect 19700 11940 19724 11942
rect 19780 11940 19786 11942
rect 19478 11920 19786 11940
rect 19478 10908 19786 10928
rect 19478 10906 19484 10908
rect 19540 10906 19564 10908
rect 19620 10906 19644 10908
rect 19700 10906 19724 10908
rect 19780 10906 19786 10908
rect 19540 10854 19542 10906
rect 19722 10854 19724 10906
rect 19478 10852 19484 10854
rect 19540 10852 19564 10854
rect 19620 10852 19644 10854
rect 19700 10852 19724 10854
rect 19780 10852 19786 10854
rect 19478 10832 19786 10852
rect 19904 10674 19932 12106
rect 19996 11762 20024 12174
rect 19984 11756 20036 11762
rect 19984 11698 20036 11704
rect 20088 11082 20116 12718
rect 20076 11076 20128 11082
rect 20076 11018 20128 11024
rect 19892 10668 19944 10674
rect 19892 10610 19944 10616
rect 20076 10668 20128 10674
rect 20076 10610 20128 10616
rect 19352 10538 19472 10554
rect 19352 10532 19484 10538
rect 19352 10526 19432 10532
rect 19432 10474 19484 10480
rect 19340 10464 19392 10470
rect 19340 10406 19392 10412
rect 19248 10124 19300 10130
rect 19248 10066 19300 10072
rect 19352 10062 19380 10406
rect 19156 10056 19208 10062
rect 19156 9998 19208 10004
rect 19340 10056 19392 10062
rect 19340 9998 19392 10004
rect 19478 9820 19786 9840
rect 19478 9818 19484 9820
rect 19540 9818 19564 9820
rect 19620 9818 19644 9820
rect 19700 9818 19724 9820
rect 19780 9818 19786 9820
rect 19540 9766 19542 9818
rect 19722 9766 19724 9818
rect 19478 9764 19484 9766
rect 19540 9764 19564 9766
rect 19620 9764 19644 9766
rect 19700 9764 19724 9766
rect 19780 9764 19786 9766
rect 19478 9744 19786 9764
rect 20088 9722 20116 10610
rect 18616 9646 18736 9674
rect 20076 9716 20128 9722
rect 20076 9658 20128 9664
rect 18052 8084 18104 8090
rect 18052 8026 18104 8032
rect 18328 8084 18380 8090
rect 18328 8026 18380 8032
rect 18512 8084 18564 8090
rect 18512 8026 18564 8032
rect 17960 6452 18012 6458
rect 17960 6394 18012 6400
rect 18064 6390 18092 8026
rect 18340 7886 18368 8026
rect 18328 7880 18380 7886
rect 18328 7822 18380 7828
rect 18524 7750 18552 8026
rect 18616 8022 18644 9646
rect 19708 9376 19760 9382
rect 19708 9318 19760 9324
rect 19720 9042 19748 9318
rect 19708 9036 19760 9042
rect 19708 8978 19760 8984
rect 19892 8968 19944 8974
rect 19892 8910 19944 8916
rect 19478 8732 19786 8752
rect 19478 8730 19484 8732
rect 19540 8730 19564 8732
rect 19620 8730 19644 8732
rect 19700 8730 19724 8732
rect 19780 8730 19786 8732
rect 19540 8678 19542 8730
rect 19722 8678 19724 8730
rect 19478 8676 19484 8678
rect 19540 8676 19564 8678
rect 19620 8676 19644 8678
rect 19700 8676 19724 8678
rect 19780 8676 19786 8678
rect 19478 8656 19786 8676
rect 19904 8566 19932 8910
rect 20076 8628 20128 8634
rect 20076 8570 20128 8576
rect 19156 8560 19208 8566
rect 19156 8502 19208 8508
rect 19432 8560 19484 8566
rect 19432 8502 19484 8508
rect 19892 8560 19944 8566
rect 19892 8502 19944 8508
rect 18694 8392 18750 8401
rect 18694 8327 18696 8336
rect 18748 8327 18750 8336
rect 18696 8298 18748 8304
rect 18604 8016 18656 8022
rect 18604 7958 18656 7964
rect 19168 7954 19196 8502
rect 19340 8356 19392 8362
rect 19340 8298 19392 8304
rect 19352 7954 19380 8298
rect 19156 7948 19208 7954
rect 19156 7890 19208 7896
rect 19340 7948 19392 7954
rect 19340 7890 19392 7896
rect 18512 7744 18564 7750
rect 19444 7732 19472 8502
rect 19984 8492 20036 8498
rect 19984 8434 20036 8440
rect 19892 8288 19944 8294
rect 19892 8230 19944 8236
rect 19616 8016 19668 8022
rect 19616 7958 19668 7964
rect 19628 7886 19656 7958
rect 19616 7880 19668 7886
rect 19616 7822 19668 7828
rect 18512 7686 18564 7692
rect 19352 7704 19472 7732
rect 18420 7200 18472 7206
rect 18420 7142 18472 7148
rect 18432 7002 18460 7142
rect 18420 6996 18472 7002
rect 18420 6938 18472 6944
rect 18052 6384 18104 6390
rect 18052 6326 18104 6332
rect 17776 6248 17828 6254
rect 17776 6190 17828 6196
rect 17788 5778 17816 6190
rect 17868 6112 17920 6118
rect 17868 6054 17920 6060
rect 17776 5772 17828 5778
rect 17776 5714 17828 5720
rect 17880 5710 17908 6054
rect 18064 5794 18092 6326
rect 17972 5766 18092 5794
rect 17972 5710 18000 5766
rect 17868 5704 17920 5710
rect 17868 5646 17920 5652
rect 17960 5704 18012 5710
rect 17960 5646 18012 5652
rect 18328 5704 18380 5710
rect 18328 5646 18380 5652
rect 18144 5636 18196 5642
rect 18144 5578 18196 5584
rect 17868 5568 17920 5574
rect 17868 5510 17920 5516
rect 17880 5370 17908 5510
rect 17868 5364 17920 5370
rect 17868 5306 17920 5312
rect 17592 5296 17644 5302
rect 17592 5238 17644 5244
rect 17960 5024 18012 5030
rect 17960 4966 18012 4972
rect 17408 4820 17460 4826
rect 17408 4762 17460 4768
rect 17224 4616 17276 4622
rect 17224 4558 17276 4564
rect 17236 4146 17264 4558
rect 17420 4146 17448 4762
rect 17776 4548 17828 4554
rect 17776 4490 17828 4496
rect 17788 4146 17816 4490
rect 17224 4140 17276 4146
rect 17224 4082 17276 4088
rect 17408 4140 17460 4146
rect 17408 4082 17460 4088
rect 17776 4140 17828 4146
rect 17776 4082 17828 4088
rect 17420 3398 17448 4082
rect 17788 3738 17816 4082
rect 17776 3732 17828 3738
rect 17776 3674 17828 3680
rect 17972 3534 18000 4966
rect 18156 4826 18184 5578
rect 18340 5370 18368 5646
rect 18328 5364 18380 5370
rect 18328 5306 18380 5312
rect 18340 5234 18368 5306
rect 18328 5228 18380 5234
rect 18328 5170 18380 5176
rect 18144 4820 18196 4826
rect 18144 4762 18196 4768
rect 18420 4616 18472 4622
rect 18420 4558 18472 4564
rect 18144 4548 18196 4554
rect 18144 4490 18196 4496
rect 18156 4146 18184 4490
rect 18144 4140 18196 4146
rect 18144 4082 18196 4088
rect 18156 3534 18184 4082
rect 18432 3738 18460 4558
rect 18420 3732 18472 3738
rect 18420 3674 18472 3680
rect 17960 3528 18012 3534
rect 17960 3470 18012 3476
rect 18144 3528 18196 3534
rect 18144 3470 18196 3476
rect 17408 3392 17460 3398
rect 17408 3334 17460 3340
rect 17052 2746 17172 2774
rect 17052 2650 17080 2746
rect 17040 2644 17092 2650
rect 17040 2586 17092 2592
rect 18524 2514 18552 7686
rect 19352 7410 19380 7704
rect 19478 7644 19786 7664
rect 19478 7642 19484 7644
rect 19540 7642 19564 7644
rect 19620 7642 19644 7644
rect 19700 7642 19724 7644
rect 19780 7642 19786 7644
rect 19540 7590 19542 7642
rect 19722 7590 19724 7642
rect 19478 7588 19484 7590
rect 19540 7588 19564 7590
rect 19620 7588 19644 7590
rect 19700 7588 19724 7590
rect 19780 7588 19786 7590
rect 19478 7568 19786 7588
rect 19340 7404 19392 7410
rect 19340 7346 19392 7352
rect 19708 7404 19760 7410
rect 19708 7346 19760 7352
rect 19064 7200 19116 7206
rect 19064 7142 19116 7148
rect 18696 6792 18748 6798
rect 18696 6734 18748 6740
rect 18708 6458 18736 6734
rect 18696 6452 18748 6458
rect 18696 6394 18748 6400
rect 18604 6384 18656 6390
rect 18604 6326 18656 6332
rect 18616 5234 18644 6326
rect 18972 6316 19024 6322
rect 18972 6258 19024 6264
rect 18788 5840 18840 5846
rect 18788 5782 18840 5788
rect 18604 5228 18656 5234
rect 18604 5170 18656 5176
rect 18616 4078 18644 5170
rect 18800 4554 18828 5782
rect 18984 5574 19012 6258
rect 19076 6118 19104 7142
rect 19248 6792 19300 6798
rect 19248 6734 19300 6740
rect 19524 6792 19576 6798
rect 19524 6734 19576 6740
rect 19064 6112 19116 6118
rect 19064 6054 19116 6060
rect 19076 5914 19104 6054
rect 19064 5908 19116 5914
rect 19064 5850 19116 5856
rect 18972 5568 19024 5574
rect 18972 5510 19024 5516
rect 18984 4622 19012 5510
rect 19260 5234 19288 6734
rect 19536 6644 19564 6734
rect 19720 6730 19748 7346
rect 19708 6724 19760 6730
rect 19708 6666 19760 6672
rect 19398 6616 19564 6644
rect 19398 6610 19426 6616
rect 19352 6582 19426 6610
rect 19352 5642 19380 6582
rect 19478 6556 19786 6576
rect 19478 6554 19484 6556
rect 19540 6554 19564 6556
rect 19620 6554 19644 6556
rect 19700 6554 19724 6556
rect 19780 6554 19786 6556
rect 19540 6502 19542 6554
rect 19722 6502 19724 6554
rect 19478 6500 19484 6502
rect 19540 6500 19564 6502
rect 19620 6500 19644 6502
rect 19700 6500 19724 6502
rect 19780 6500 19786 6502
rect 19478 6480 19786 6500
rect 19432 6180 19484 6186
rect 19432 6122 19484 6128
rect 19444 5914 19472 6122
rect 19432 5908 19484 5914
rect 19432 5850 19484 5856
rect 19904 5778 19932 8230
rect 19996 8090 20024 8434
rect 19984 8084 20036 8090
rect 19984 8026 20036 8032
rect 19984 7880 20036 7886
rect 19984 7822 20036 7828
rect 19996 7478 20024 7822
rect 19984 7472 20036 7478
rect 19984 7414 20036 7420
rect 19984 7336 20036 7342
rect 19984 7278 20036 7284
rect 19996 6662 20024 7278
rect 19984 6656 20036 6662
rect 19984 6598 20036 6604
rect 19996 6322 20024 6598
rect 19984 6316 20036 6322
rect 19984 6258 20036 6264
rect 20088 6186 20116 8570
rect 20076 6180 20128 6186
rect 20076 6122 20128 6128
rect 19892 5772 19944 5778
rect 19892 5714 19944 5720
rect 19340 5636 19392 5642
rect 19340 5578 19392 5584
rect 19478 5468 19786 5488
rect 19478 5466 19484 5468
rect 19540 5466 19564 5468
rect 19620 5466 19644 5468
rect 19700 5466 19724 5468
rect 19780 5466 19786 5468
rect 19540 5414 19542 5466
rect 19722 5414 19724 5466
rect 19478 5412 19484 5414
rect 19540 5412 19564 5414
rect 19620 5412 19644 5414
rect 19700 5412 19724 5414
rect 19780 5412 19786 5414
rect 19478 5392 19786 5412
rect 19904 5370 19932 5714
rect 19892 5364 19944 5370
rect 19892 5306 19944 5312
rect 19248 5228 19300 5234
rect 19248 5170 19300 5176
rect 19260 5030 19288 5170
rect 19248 5024 19300 5030
rect 19248 4966 19300 4972
rect 18972 4616 19024 4622
rect 18972 4558 19024 4564
rect 18788 4548 18840 4554
rect 18788 4490 18840 4496
rect 18984 4214 19012 4558
rect 19340 4480 19392 4486
rect 19340 4422 19392 4428
rect 19352 4282 19380 4422
rect 19478 4380 19786 4400
rect 19478 4378 19484 4380
rect 19540 4378 19564 4380
rect 19620 4378 19644 4380
rect 19700 4378 19724 4380
rect 19780 4378 19786 4380
rect 19540 4326 19542 4378
rect 19722 4326 19724 4378
rect 19478 4324 19484 4326
rect 19540 4324 19564 4326
rect 19620 4324 19644 4326
rect 19700 4324 19724 4326
rect 19780 4324 19786 4326
rect 19478 4304 19786 4324
rect 19340 4276 19392 4282
rect 19340 4218 19392 4224
rect 18972 4208 19024 4214
rect 18972 4150 19024 4156
rect 18604 4072 18656 4078
rect 18604 4014 18656 4020
rect 18616 3602 18644 4014
rect 18984 3738 19012 4150
rect 19904 4146 19932 5306
rect 19984 4548 20036 4554
rect 19984 4490 20036 4496
rect 19708 4140 19760 4146
rect 19708 4082 19760 4088
rect 19892 4140 19944 4146
rect 19892 4082 19944 4088
rect 19248 3936 19300 3942
rect 19248 3878 19300 3884
rect 18972 3732 19024 3738
rect 18972 3674 19024 3680
rect 19260 3670 19288 3878
rect 19248 3664 19300 3670
rect 19248 3606 19300 3612
rect 18604 3596 18656 3602
rect 18604 3538 18656 3544
rect 19260 3534 19288 3606
rect 19720 3534 19748 4082
rect 19904 3602 19932 4082
rect 19892 3596 19944 3602
rect 19892 3538 19944 3544
rect 19248 3528 19300 3534
rect 19248 3470 19300 3476
rect 19708 3528 19760 3534
rect 19708 3470 19760 3476
rect 19478 3292 19786 3312
rect 19478 3290 19484 3292
rect 19540 3290 19564 3292
rect 19620 3290 19644 3292
rect 19700 3290 19724 3292
rect 19780 3290 19786 3292
rect 19540 3238 19542 3290
rect 19722 3238 19724 3290
rect 19478 3236 19484 3238
rect 19540 3236 19564 3238
rect 19620 3236 19644 3238
rect 19700 3236 19724 3238
rect 19780 3236 19786 3238
rect 19478 3216 19786 3236
rect 19904 3126 19932 3538
rect 19996 3398 20024 4490
rect 20076 4480 20128 4486
rect 20076 4422 20128 4428
rect 19984 3392 20036 3398
rect 19984 3334 20036 3340
rect 19892 3120 19944 3126
rect 19892 3062 19944 3068
rect 20088 3058 20116 4422
rect 20076 3052 20128 3058
rect 20076 2994 20128 3000
rect 20180 2774 20208 12786
rect 20272 11778 20300 16594
rect 20352 16040 20404 16046
rect 20352 15982 20404 15988
rect 20364 15570 20392 15982
rect 20352 15564 20404 15570
rect 20352 15506 20404 15512
rect 20456 15201 20484 16918
rect 20732 16522 20760 16934
rect 21100 16590 21128 17274
rect 21192 17202 21220 18702
rect 21732 18692 21784 18698
rect 21732 18634 21784 18640
rect 21640 17876 21692 17882
rect 21640 17818 21692 17824
rect 21272 17672 21324 17678
rect 21272 17614 21324 17620
rect 21180 17196 21232 17202
rect 21180 17138 21232 17144
rect 21088 16584 21140 16590
rect 21088 16526 21140 16532
rect 20720 16516 20772 16522
rect 20720 16458 20772 16464
rect 21180 16516 21232 16522
rect 21180 16458 21232 16464
rect 21088 16448 21140 16454
rect 21088 16390 21140 16396
rect 20994 16144 21050 16153
rect 21100 16114 21128 16390
rect 21192 16250 21220 16458
rect 21180 16244 21232 16250
rect 21180 16186 21232 16192
rect 20994 16079 21050 16088
rect 21088 16108 21140 16114
rect 21008 15978 21036 16079
rect 21088 16050 21140 16056
rect 20996 15972 21048 15978
rect 20996 15914 21048 15920
rect 21088 15972 21140 15978
rect 21088 15914 21140 15920
rect 21100 15858 21128 15914
rect 20916 15830 21128 15858
rect 20536 15632 20588 15638
rect 20536 15574 20588 15580
rect 20442 15192 20498 15201
rect 20442 15127 20444 15136
rect 20496 15127 20498 15136
rect 20444 15098 20496 15104
rect 20456 15067 20484 15098
rect 20548 14958 20576 15574
rect 20720 15428 20772 15434
rect 20720 15370 20772 15376
rect 20628 15088 20680 15094
rect 20732 15065 20760 15370
rect 20628 15030 20680 15036
rect 20718 15056 20774 15065
rect 20536 14952 20588 14958
rect 20536 14894 20588 14900
rect 20548 14550 20576 14894
rect 20640 14550 20668 15030
rect 20718 14991 20720 15000
rect 20772 14991 20774 15000
rect 20720 14962 20772 14968
rect 20536 14544 20588 14550
rect 20536 14486 20588 14492
rect 20628 14544 20680 14550
rect 20628 14486 20680 14492
rect 20536 14340 20588 14346
rect 20536 14282 20588 14288
rect 20352 14272 20404 14278
rect 20352 14214 20404 14220
rect 20364 14074 20392 14214
rect 20352 14068 20404 14074
rect 20352 14010 20404 14016
rect 20548 14006 20576 14282
rect 20732 14278 20760 14962
rect 20720 14272 20772 14278
rect 20720 14214 20772 14220
rect 20536 14000 20588 14006
rect 20536 13942 20588 13948
rect 20916 13938 20944 15830
rect 21088 15496 21140 15502
rect 21088 15438 21140 15444
rect 20996 15020 21048 15026
rect 20996 14962 21048 14968
rect 21008 14346 21036 14962
rect 21100 14890 21128 15438
rect 21284 15162 21312 17614
rect 21364 17196 21416 17202
rect 21364 17138 21416 17144
rect 21272 15156 21324 15162
rect 21272 15098 21324 15104
rect 21180 15020 21232 15026
rect 21180 14962 21232 14968
rect 21192 14890 21220 14962
rect 21088 14884 21140 14890
rect 21088 14826 21140 14832
rect 21180 14884 21232 14890
rect 21180 14826 21232 14832
rect 21192 14414 21220 14826
rect 21376 14618 21404 17138
rect 21548 15904 21600 15910
rect 21548 15846 21600 15852
rect 21456 15564 21508 15570
rect 21456 15506 21508 15512
rect 21364 14612 21416 14618
rect 21364 14554 21416 14560
rect 21468 14482 21496 15506
rect 21456 14476 21508 14482
rect 21456 14418 21508 14424
rect 21180 14408 21232 14414
rect 21180 14350 21232 14356
rect 20996 14340 21048 14346
rect 20996 14282 21048 14288
rect 21192 13938 21220 14350
rect 20904 13932 20956 13938
rect 20904 13874 20956 13880
rect 21180 13932 21232 13938
rect 21180 13874 21232 13880
rect 20536 13524 20588 13530
rect 20536 13466 20588 13472
rect 20352 13252 20404 13258
rect 20352 13194 20404 13200
rect 20364 12442 20392 13194
rect 20444 12980 20496 12986
rect 20444 12922 20496 12928
rect 20352 12436 20404 12442
rect 20352 12378 20404 12384
rect 20456 11898 20484 12922
rect 20548 12434 20576 13466
rect 20916 13462 20944 13874
rect 20904 13456 20956 13462
rect 20904 13398 20956 13404
rect 21192 13326 21220 13874
rect 21180 13320 21232 13326
rect 21180 13262 21232 13268
rect 20720 13184 20772 13190
rect 20720 13126 20772 13132
rect 21180 13184 21232 13190
rect 21180 13126 21232 13132
rect 20548 12406 20668 12434
rect 20444 11892 20496 11898
rect 20444 11834 20496 11840
rect 20272 11750 20392 11778
rect 20260 11688 20312 11694
rect 20260 11630 20312 11636
rect 20364 11642 20392 11750
rect 20272 10810 20300 11630
rect 20364 11614 20484 11642
rect 20352 11552 20404 11558
rect 20352 11494 20404 11500
rect 20260 10804 20312 10810
rect 20260 10746 20312 10752
rect 20364 10674 20392 11494
rect 20352 10668 20404 10674
rect 20352 10610 20404 10616
rect 20352 10532 20404 10538
rect 20352 10474 20404 10480
rect 20260 7744 20312 7750
rect 20260 7686 20312 7692
rect 20272 6390 20300 7686
rect 20364 6746 20392 10474
rect 20456 8906 20484 11614
rect 20536 11620 20588 11626
rect 20536 11562 20588 11568
rect 20548 9518 20576 11562
rect 20536 9512 20588 9518
rect 20536 9454 20588 9460
rect 20444 8900 20496 8906
rect 20444 8842 20496 8848
rect 20536 8832 20588 8838
rect 20536 8774 20588 8780
rect 20548 8022 20576 8774
rect 20640 8090 20668 12406
rect 20732 11762 20760 13126
rect 20904 12912 20956 12918
rect 20904 12854 20956 12860
rect 20810 12336 20866 12345
rect 20810 12271 20866 12280
rect 20824 12238 20852 12271
rect 20812 12232 20864 12238
rect 20812 12174 20864 12180
rect 20916 12084 20944 12854
rect 21192 12850 21220 13126
rect 21088 12844 21140 12850
rect 21088 12786 21140 12792
rect 21180 12844 21232 12850
rect 21180 12786 21232 12792
rect 20824 12056 20944 12084
rect 20720 11756 20772 11762
rect 20720 11698 20772 11704
rect 20824 11354 20852 12056
rect 21100 11898 21128 12786
rect 21192 12306 21220 12786
rect 21456 12640 21508 12646
rect 21456 12582 21508 12588
rect 21180 12300 21232 12306
rect 21180 12242 21232 12248
rect 20904 11892 20956 11898
rect 20904 11834 20956 11840
rect 21088 11892 21140 11898
rect 21088 11834 21140 11840
rect 20812 11348 20864 11354
rect 20812 11290 20864 11296
rect 20916 10674 20944 11834
rect 20996 11824 21048 11830
rect 20996 11766 21048 11772
rect 21008 11354 21036 11766
rect 21192 11694 21220 12242
rect 21364 12232 21416 12238
rect 21364 12174 21416 12180
rect 21180 11688 21232 11694
rect 21180 11630 21232 11636
rect 21180 11552 21232 11558
rect 21180 11494 21232 11500
rect 20996 11348 21048 11354
rect 20996 11290 21048 11296
rect 21008 10810 21036 11290
rect 20996 10804 21048 10810
rect 20996 10746 21048 10752
rect 21192 10742 21220 11494
rect 21376 10742 21404 12174
rect 21468 12102 21496 12582
rect 21456 12096 21508 12102
rect 21456 12038 21508 12044
rect 21180 10736 21232 10742
rect 21180 10678 21232 10684
rect 21364 10736 21416 10742
rect 21364 10678 21416 10684
rect 21468 10674 21496 12038
rect 20904 10668 20956 10674
rect 20904 10610 20956 10616
rect 21456 10668 21508 10674
rect 21456 10610 21508 10616
rect 21180 9920 21232 9926
rect 21180 9862 21232 9868
rect 21192 9654 21220 9862
rect 21180 9648 21232 9654
rect 21180 9590 21232 9596
rect 21272 9580 21324 9586
rect 21272 9522 21324 9528
rect 21284 9178 21312 9522
rect 21272 9172 21324 9178
rect 21272 9114 21324 9120
rect 20996 9104 21048 9110
rect 20996 9046 21048 9052
rect 20720 8968 20772 8974
rect 20720 8910 20772 8916
rect 20732 8634 20760 8910
rect 20720 8628 20772 8634
rect 20720 8570 20772 8576
rect 20628 8084 20680 8090
rect 20628 8026 20680 8032
rect 20536 8016 20588 8022
rect 20536 7958 20588 7964
rect 20548 7886 20576 7958
rect 21008 7886 21036 9046
rect 21088 8356 21140 8362
rect 21088 8298 21140 8304
rect 20444 7880 20496 7886
rect 20444 7822 20496 7828
rect 20536 7880 20588 7886
rect 20536 7822 20588 7828
rect 20996 7880 21048 7886
rect 20996 7822 21048 7828
rect 20456 6866 20484 7822
rect 20628 7812 20680 7818
rect 20628 7754 20680 7760
rect 20640 7698 20668 7754
rect 20904 7744 20956 7750
rect 20640 7670 20760 7698
rect 20904 7686 20956 7692
rect 20536 7472 20588 7478
rect 20536 7414 20588 7420
rect 20548 7002 20576 7414
rect 20536 6996 20588 7002
rect 20536 6938 20588 6944
rect 20444 6860 20496 6866
rect 20444 6802 20496 6808
rect 20364 6718 20484 6746
rect 20260 6384 20312 6390
rect 20260 6326 20312 6332
rect 20272 6202 20300 6326
rect 20272 6174 20392 6202
rect 20260 6112 20312 6118
rect 20260 6054 20312 6060
rect 20272 5710 20300 6054
rect 20260 5704 20312 5710
rect 20260 5646 20312 5652
rect 20364 5574 20392 6174
rect 20352 5568 20404 5574
rect 20352 5510 20404 5516
rect 20364 4622 20392 5510
rect 20352 4616 20404 4622
rect 20352 4558 20404 4564
rect 20352 3460 20404 3466
rect 20352 3402 20404 3408
rect 20364 3194 20392 3402
rect 20352 3188 20404 3194
rect 20352 3130 20404 3136
rect 20180 2746 20392 2774
rect 20364 2514 20392 2746
rect 20456 2582 20484 6718
rect 20548 4826 20576 6938
rect 20536 4820 20588 4826
rect 20536 4762 20588 4768
rect 20548 4622 20576 4762
rect 20536 4616 20588 4622
rect 20536 4558 20588 4564
rect 20628 4480 20680 4486
rect 20628 4422 20680 4428
rect 20640 4214 20668 4422
rect 20628 4208 20680 4214
rect 20628 4150 20680 4156
rect 20732 2650 20760 7670
rect 20916 7546 20944 7686
rect 20904 7540 20956 7546
rect 20904 7482 20956 7488
rect 21008 7478 21036 7822
rect 20996 7472 21048 7478
rect 20996 7414 21048 7420
rect 20812 7404 20864 7410
rect 20812 7346 20864 7352
rect 20824 6798 20852 7346
rect 21100 6798 21128 8298
rect 21560 7970 21588 15846
rect 21652 15178 21680 17818
rect 21744 17610 21772 18634
rect 21836 18630 21864 18838
rect 22284 18760 22336 18766
rect 22284 18702 22336 18708
rect 21824 18624 21876 18630
rect 21824 18566 21876 18572
rect 22008 18624 22060 18630
rect 22008 18566 22060 18572
rect 21916 18352 21968 18358
rect 21916 18294 21968 18300
rect 21824 18284 21876 18290
rect 21824 18226 21876 18232
rect 21732 17604 21784 17610
rect 21732 17546 21784 17552
rect 21744 16998 21772 17546
rect 21732 16992 21784 16998
rect 21732 16934 21784 16940
rect 21732 16584 21784 16590
rect 21836 16572 21864 18226
rect 21928 17542 21956 18294
rect 22020 18290 22048 18566
rect 22100 18420 22152 18426
rect 22100 18362 22152 18368
rect 22008 18284 22060 18290
rect 22008 18226 22060 18232
rect 22112 17649 22140 18362
rect 22296 18290 22324 18702
rect 22480 18426 22508 20810
rect 22744 20052 22796 20058
rect 22744 19994 22796 20000
rect 22652 19780 22704 19786
rect 22652 19722 22704 19728
rect 22664 19514 22692 19722
rect 22652 19508 22704 19514
rect 22652 19450 22704 19456
rect 22652 19304 22704 19310
rect 22652 19246 22704 19252
rect 22664 18630 22692 19246
rect 22652 18624 22704 18630
rect 22652 18566 22704 18572
rect 22468 18420 22520 18426
rect 22468 18362 22520 18368
rect 22284 18284 22336 18290
rect 22284 18226 22336 18232
rect 22296 17814 22324 18226
rect 22664 18154 22692 18566
rect 22756 18358 22784 19994
rect 22744 18352 22796 18358
rect 22744 18294 22796 18300
rect 22652 18148 22704 18154
rect 22652 18090 22704 18096
rect 22284 17808 22336 17814
rect 22284 17750 22336 17756
rect 22098 17640 22154 17649
rect 22098 17575 22154 17584
rect 22468 17604 22520 17610
rect 22468 17546 22520 17552
rect 21916 17536 21968 17542
rect 21916 17478 21968 17484
rect 22192 17196 22244 17202
rect 22192 17138 22244 17144
rect 21916 16992 21968 16998
rect 21916 16934 21968 16940
rect 21928 16590 21956 16934
rect 21784 16544 21864 16572
rect 21916 16584 21968 16590
rect 21732 16526 21784 16532
rect 21916 16526 21968 16532
rect 21744 16114 21772 16526
rect 22204 16522 22232 17138
rect 22480 16590 22508 17546
rect 22664 16726 22692 18090
rect 22756 17746 22784 18294
rect 22744 17740 22796 17746
rect 22744 17682 22796 17688
rect 22652 16720 22704 16726
rect 22652 16662 22704 16668
rect 22468 16584 22520 16590
rect 22468 16526 22520 16532
rect 22192 16516 22244 16522
rect 22192 16458 22244 16464
rect 22480 16182 22508 16526
rect 22560 16516 22612 16522
rect 22560 16458 22612 16464
rect 22468 16176 22520 16182
rect 22468 16118 22520 16124
rect 21732 16108 21784 16114
rect 21732 16050 21784 16056
rect 22008 16108 22060 16114
rect 22008 16050 22060 16056
rect 22020 15706 22048 16050
rect 22098 16008 22154 16017
rect 22098 15943 22100 15952
rect 22152 15943 22154 15952
rect 22100 15914 22152 15920
rect 22008 15700 22060 15706
rect 22008 15642 22060 15648
rect 22192 15700 22244 15706
rect 22192 15642 22244 15648
rect 22006 15464 22062 15473
rect 21916 15428 21968 15434
rect 22006 15399 22062 15408
rect 21916 15370 21968 15376
rect 21652 15150 21864 15178
rect 21732 15020 21784 15026
rect 21732 14962 21784 14968
rect 21640 14408 21692 14414
rect 21640 14350 21692 14356
rect 21652 13190 21680 14350
rect 21744 13734 21772 14962
rect 21732 13728 21784 13734
rect 21732 13670 21784 13676
rect 21744 13326 21772 13670
rect 21732 13320 21784 13326
rect 21732 13262 21784 13268
rect 21640 13184 21692 13190
rect 21640 13126 21692 13132
rect 21652 12238 21680 13126
rect 21836 12442 21864 15150
rect 21928 15094 21956 15370
rect 22020 15314 22048 15399
rect 22020 15286 22140 15314
rect 22008 15156 22060 15162
rect 22008 15098 22060 15104
rect 21916 15088 21968 15094
rect 21916 15030 21968 15036
rect 22020 14958 22048 15098
rect 22008 14952 22060 14958
rect 22008 14894 22060 14900
rect 22008 14408 22060 14414
rect 22008 14350 22060 14356
rect 22020 13530 22048 14350
rect 22008 13524 22060 13530
rect 22008 13466 22060 13472
rect 21824 12436 21876 12442
rect 21824 12378 21876 12384
rect 21640 12232 21692 12238
rect 21640 12174 21692 12180
rect 21916 12096 21968 12102
rect 21916 12038 21968 12044
rect 21928 11830 21956 12038
rect 21916 11824 21968 11830
rect 21916 11766 21968 11772
rect 22112 11762 22140 15286
rect 22204 12306 22232 15642
rect 22480 15638 22508 16118
rect 22468 15632 22520 15638
rect 22468 15574 22520 15580
rect 22376 15496 22428 15502
rect 22376 15438 22428 15444
rect 22388 14346 22416 15438
rect 22572 15366 22600 16458
rect 22652 15496 22704 15502
rect 22652 15438 22704 15444
rect 22560 15360 22612 15366
rect 22560 15302 22612 15308
rect 22572 14618 22600 15302
rect 22560 14612 22612 14618
rect 22560 14554 22612 14560
rect 22664 14414 22692 15438
rect 22652 14408 22704 14414
rect 22652 14350 22704 14356
rect 22376 14340 22428 14346
rect 22376 14282 22428 14288
rect 22560 13728 22612 13734
rect 22560 13670 22612 13676
rect 22284 13388 22336 13394
rect 22284 13330 22336 13336
rect 22296 12714 22324 13330
rect 22468 13320 22520 13326
rect 22466 13288 22468 13297
rect 22520 13288 22522 13297
rect 22466 13223 22522 13232
rect 22572 13172 22600 13670
rect 22652 13184 22704 13190
rect 22572 13144 22652 13172
rect 22652 13126 22704 13132
rect 22284 12708 22336 12714
rect 22284 12650 22336 12656
rect 22296 12306 22324 12650
rect 22192 12300 22244 12306
rect 22192 12242 22244 12248
rect 22284 12300 22336 12306
rect 22284 12242 22336 12248
rect 22558 12200 22614 12209
rect 22558 12135 22560 12144
rect 22612 12135 22614 12144
rect 22560 12106 22612 12112
rect 22100 11756 22152 11762
rect 22100 11698 22152 11704
rect 22376 11756 22428 11762
rect 22376 11698 22428 11704
rect 22112 11354 22140 11698
rect 22100 11348 22152 11354
rect 22100 11290 22152 11296
rect 21916 10464 21968 10470
rect 21916 10406 21968 10412
rect 21928 10130 21956 10406
rect 21916 10124 21968 10130
rect 21916 10066 21968 10072
rect 22008 9920 22060 9926
rect 22008 9862 22060 9868
rect 22020 9722 22048 9862
rect 22008 9716 22060 9722
rect 22008 9658 22060 9664
rect 21732 9104 21784 9110
rect 21732 9046 21784 9052
rect 21640 8968 21692 8974
rect 21640 8910 21692 8916
rect 21652 8634 21680 8910
rect 21640 8628 21692 8634
rect 21640 8570 21692 8576
rect 21744 8022 21772 9046
rect 22020 8974 22048 9658
rect 22008 8968 22060 8974
rect 22008 8910 22060 8916
rect 21824 8832 21876 8838
rect 21824 8774 21876 8780
rect 21468 7942 21588 7970
rect 21732 8016 21784 8022
rect 21732 7958 21784 7964
rect 21180 7744 21232 7750
rect 21364 7744 21416 7750
rect 21232 7692 21364 7698
rect 21180 7686 21416 7692
rect 21192 7670 21404 7686
rect 21180 7472 21232 7478
rect 21180 7414 21232 7420
rect 20812 6792 20864 6798
rect 20812 6734 20864 6740
rect 21088 6792 21140 6798
rect 21088 6734 21140 6740
rect 21100 6322 21128 6734
rect 21088 6316 21140 6322
rect 21088 6258 21140 6264
rect 20996 6180 21048 6186
rect 20996 6122 21048 6128
rect 21008 5778 21036 6122
rect 20996 5772 21048 5778
rect 20996 5714 21048 5720
rect 21192 4690 21220 7414
rect 21376 7274 21404 7670
rect 21364 7268 21416 7274
rect 21364 7210 21416 7216
rect 21272 6792 21324 6798
rect 21272 6734 21324 6740
rect 21284 6458 21312 6734
rect 21272 6452 21324 6458
rect 21272 6394 21324 6400
rect 21284 5914 21312 6394
rect 21376 6254 21404 7210
rect 21364 6248 21416 6254
rect 21364 6190 21416 6196
rect 21272 5908 21324 5914
rect 21272 5850 21324 5856
rect 21376 5710 21404 6190
rect 21364 5704 21416 5710
rect 21364 5646 21416 5652
rect 21180 4684 21232 4690
rect 21180 4626 21232 4632
rect 21468 3534 21496 7942
rect 21640 7336 21692 7342
rect 21640 7278 21692 7284
rect 21652 6730 21680 7278
rect 21744 7206 21772 7958
rect 21836 7478 21864 8774
rect 21824 7472 21876 7478
rect 21824 7414 21876 7420
rect 21732 7200 21784 7206
rect 21732 7142 21784 7148
rect 22112 6866 22140 11290
rect 22388 10266 22416 11698
rect 22560 11552 22612 11558
rect 22560 11494 22612 11500
rect 22572 11082 22600 11494
rect 22560 11076 22612 11082
rect 22560 11018 22612 11024
rect 22468 11008 22520 11014
rect 22468 10950 22520 10956
rect 22480 10742 22508 10950
rect 22468 10736 22520 10742
rect 22468 10678 22520 10684
rect 22560 10600 22612 10606
rect 22560 10542 22612 10548
rect 22572 10266 22600 10542
rect 22376 10260 22428 10266
rect 22376 10202 22428 10208
rect 22560 10260 22612 10266
rect 22560 10202 22612 10208
rect 22468 10056 22520 10062
rect 22468 9998 22520 10004
rect 22480 9722 22508 9998
rect 22468 9716 22520 9722
rect 22468 9658 22520 9664
rect 22572 9654 22600 10202
rect 22560 9648 22612 9654
rect 22560 9590 22612 9596
rect 22192 9580 22244 9586
rect 22192 9522 22244 9528
rect 22204 9178 22232 9522
rect 22192 9172 22244 9178
rect 22192 9114 22244 9120
rect 22664 8566 22692 13126
rect 22756 12986 22784 17682
rect 22848 15994 22876 23802
rect 23952 22094 23980 26206
rect 24110 25596 24418 25616
rect 24110 25594 24116 25596
rect 24172 25594 24196 25596
rect 24252 25594 24276 25596
rect 24332 25594 24356 25596
rect 24412 25594 24418 25596
rect 24172 25542 24174 25594
rect 24354 25542 24356 25594
rect 24110 25540 24116 25542
rect 24172 25540 24196 25542
rect 24252 25540 24276 25542
rect 24332 25540 24356 25542
rect 24412 25540 24418 25542
rect 24110 25520 24418 25540
rect 24110 24508 24418 24528
rect 24110 24506 24116 24508
rect 24172 24506 24196 24508
rect 24252 24506 24276 24508
rect 24332 24506 24356 24508
rect 24412 24506 24418 24508
rect 24172 24454 24174 24506
rect 24354 24454 24356 24506
rect 24110 24452 24116 24454
rect 24172 24452 24196 24454
rect 24252 24452 24276 24454
rect 24332 24452 24356 24454
rect 24412 24452 24418 24454
rect 24110 24432 24418 24452
rect 24110 23420 24418 23440
rect 24110 23418 24116 23420
rect 24172 23418 24196 23420
rect 24252 23418 24276 23420
rect 24332 23418 24356 23420
rect 24412 23418 24418 23420
rect 24172 23366 24174 23418
rect 24354 23366 24356 23418
rect 24110 23364 24116 23366
rect 24172 23364 24196 23366
rect 24252 23364 24276 23366
rect 24332 23364 24356 23366
rect 24412 23364 24418 23366
rect 24110 23344 24418 23364
rect 24110 22332 24418 22352
rect 24110 22330 24116 22332
rect 24172 22330 24196 22332
rect 24252 22330 24276 22332
rect 24332 22330 24356 22332
rect 24412 22330 24418 22332
rect 24172 22278 24174 22330
rect 24354 22278 24356 22330
rect 24110 22276 24116 22278
rect 24172 22276 24196 22278
rect 24252 22276 24276 22278
rect 24332 22276 24356 22278
rect 24412 22276 24418 22278
rect 24110 22256 24418 22276
rect 23768 22066 23980 22094
rect 23204 20936 23256 20942
rect 23204 20878 23256 20884
rect 23216 20398 23244 20878
rect 23204 20392 23256 20398
rect 23204 20334 23256 20340
rect 23020 19712 23072 19718
rect 23020 19654 23072 19660
rect 23032 19378 23060 19654
rect 23020 19372 23072 19378
rect 23020 19314 23072 19320
rect 23216 19242 23244 20334
rect 23296 19372 23348 19378
rect 23296 19314 23348 19320
rect 23664 19372 23716 19378
rect 23664 19314 23716 19320
rect 23204 19236 23256 19242
rect 23204 19178 23256 19184
rect 22928 18760 22980 18766
rect 22928 18702 22980 18708
rect 22940 18086 22968 18702
rect 23020 18284 23072 18290
rect 23020 18226 23072 18232
rect 22928 18080 22980 18086
rect 22928 18022 22980 18028
rect 22940 16572 22968 18022
rect 23032 17882 23060 18226
rect 23112 18080 23164 18086
rect 23112 18022 23164 18028
rect 23020 17876 23072 17882
rect 23020 17818 23072 17824
rect 23124 17678 23152 18022
rect 23112 17672 23164 17678
rect 23112 17614 23164 17620
rect 23020 17604 23072 17610
rect 23020 17546 23072 17552
rect 23032 17338 23060 17546
rect 23204 17536 23256 17542
rect 23308 17524 23336 19314
rect 23572 19304 23624 19310
rect 23572 19246 23624 19252
rect 23584 18766 23612 19246
rect 23676 18970 23704 19314
rect 23664 18964 23716 18970
rect 23664 18906 23716 18912
rect 23480 18760 23532 18766
rect 23480 18702 23532 18708
rect 23572 18760 23624 18766
rect 23572 18702 23624 18708
rect 23492 18630 23520 18702
rect 23480 18624 23532 18630
rect 23480 18566 23532 18572
rect 23492 18222 23520 18566
rect 23480 18216 23532 18222
rect 23480 18158 23532 18164
rect 23768 17762 23796 22066
rect 25056 21690 25084 27338
rect 25148 27130 25176 27406
rect 27540 27130 27568 29271
rect 28000 27606 28028 29294
rect 28354 29200 28410 29294
rect 29642 29200 29698 30000
rect 28262 27976 28318 27985
rect 28262 27911 28318 27920
rect 28276 27606 28304 27911
rect 27988 27600 28040 27606
rect 27988 27542 28040 27548
rect 28264 27600 28316 27606
rect 28264 27542 28316 27548
rect 25136 27124 25188 27130
rect 25136 27066 25188 27072
rect 27528 27124 27580 27130
rect 27528 27066 27580 27072
rect 28080 26988 28132 26994
rect 28080 26930 28132 26936
rect 25044 21684 25096 21690
rect 25044 21626 25096 21632
rect 24110 21244 24418 21264
rect 24110 21242 24116 21244
rect 24172 21242 24196 21244
rect 24252 21242 24276 21244
rect 24332 21242 24356 21244
rect 24412 21242 24418 21244
rect 24172 21190 24174 21242
rect 24354 21190 24356 21242
rect 24110 21188 24116 21190
rect 24172 21188 24196 21190
rect 24252 21188 24276 21190
rect 24332 21188 24356 21190
rect 24412 21188 24418 21190
rect 24110 21168 24418 21188
rect 24110 20156 24418 20176
rect 24110 20154 24116 20156
rect 24172 20154 24196 20156
rect 24252 20154 24276 20156
rect 24332 20154 24356 20156
rect 24412 20154 24418 20156
rect 24172 20102 24174 20154
rect 24354 20102 24356 20154
rect 24110 20100 24116 20102
rect 24172 20100 24196 20102
rect 24252 20100 24276 20102
rect 24332 20100 24356 20102
rect 24412 20100 24418 20102
rect 24110 20080 24418 20100
rect 24216 19848 24268 19854
rect 24216 19790 24268 19796
rect 24228 19446 24256 19790
rect 24216 19440 24268 19446
rect 24216 19382 24268 19388
rect 24676 19304 24728 19310
rect 24676 19246 24728 19252
rect 23848 19168 23900 19174
rect 23848 19110 23900 19116
rect 23940 19168 23992 19174
rect 23940 19110 23992 19116
rect 23860 18834 23888 19110
rect 23848 18828 23900 18834
rect 23848 18770 23900 18776
rect 23952 18766 23980 19110
rect 24110 19068 24418 19088
rect 24110 19066 24116 19068
rect 24172 19066 24196 19068
rect 24252 19066 24276 19068
rect 24332 19066 24356 19068
rect 24412 19066 24418 19068
rect 24172 19014 24174 19066
rect 24354 19014 24356 19066
rect 24110 19012 24116 19014
rect 24172 19012 24196 19014
rect 24252 19012 24276 19014
rect 24332 19012 24356 19014
rect 24412 19012 24418 19014
rect 24110 18992 24418 19012
rect 23940 18760 23992 18766
rect 23940 18702 23992 18708
rect 23848 18284 23900 18290
rect 23952 18272 23980 18702
rect 23900 18244 23980 18272
rect 23848 18226 23900 18232
rect 23676 17734 23796 17762
rect 23256 17496 23336 17524
rect 23388 17536 23440 17542
rect 23204 17478 23256 17484
rect 23388 17478 23440 17484
rect 23020 17332 23072 17338
rect 23020 17274 23072 17280
rect 23032 17134 23060 17274
rect 23216 17202 23244 17478
rect 23204 17196 23256 17202
rect 23204 17138 23256 17144
rect 23020 17128 23072 17134
rect 23020 17070 23072 17076
rect 23296 16652 23348 16658
rect 23216 16612 23296 16640
rect 23020 16584 23072 16590
rect 22940 16544 23020 16572
rect 23020 16526 23072 16532
rect 23032 16114 23060 16526
rect 23112 16516 23164 16522
rect 23112 16458 23164 16464
rect 23020 16108 23072 16114
rect 23020 16050 23072 16056
rect 22848 15966 22968 15994
rect 22836 15904 22888 15910
rect 22836 15846 22888 15852
rect 22744 12980 22796 12986
rect 22744 12922 22796 12928
rect 22848 12434 22876 15846
rect 22940 15706 22968 15966
rect 22928 15700 22980 15706
rect 22928 15642 22980 15648
rect 23032 15638 23060 16050
rect 23124 15978 23152 16458
rect 23216 16114 23244 16612
rect 23296 16594 23348 16600
rect 23400 16590 23428 17478
rect 23388 16584 23440 16590
rect 23572 16584 23624 16590
rect 23388 16526 23440 16532
rect 23492 16544 23572 16572
rect 23204 16108 23256 16114
rect 23388 16108 23440 16114
rect 23204 16050 23256 16056
rect 23308 16068 23388 16096
rect 23112 15972 23164 15978
rect 23112 15914 23164 15920
rect 23020 15632 23072 15638
rect 23020 15574 23072 15580
rect 23124 15620 23152 15914
rect 23204 15632 23256 15638
rect 23124 15592 23204 15620
rect 22928 15360 22980 15366
rect 22928 15302 22980 15308
rect 22940 14958 22968 15302
rect 23032 15026 23060 15574
rect 23020 15020 23072 15026
rect 23020 14962 23072 14968
rect 22928 14952 22980 14958
rect 22928 14894 22980 14900
rect 23124 14618 23152 15592
rect 23204 15574 23256 15580
rect 23112 14612 23164 14618
rect 23112 14554 23164 14560
rect 23308 13326 23336 16068
rect 23388 16050 23440 16056
rect 23492 14929 23520 16544
rect 23572 16526 23624 16532
rect 23676 16454 23704 17734
rect 23848 17604 23900 17610
rect 23768 17564 23848 17592
rect 23768 17134 23796 17564
rect 23848 17546 23900 17552
rect 23848 17196 23900 17202
rect 23848 17138 23900 17144
rect 23756 17128 23808 17134
rect 23756 17070 23808 17076
rect 23768 16522 23796 17070
rect 23860 16794 23888 17138
rect 23952 17134 23980 18244
rect 24110 17980 24418 18000
rect 24110 17978 24116 17980
rect 24172 17978 24196 17980
rect 24252 17978 24276 17980
rect 24332 17978 24356 17980
rect 24412 17978 24418 17980
rect 24172 17926 24174 17978
rect 24354 17926 24356 17978
rect 24110 17924 24116 17926
rect 24172 17924 24196 17926
rect 24252 17924 24276 17926
rect 24332 17924 24356 17926
rect 24412 17924 24418 17926
rect 24110 17904 24418 17924
rect 23940 17128 23992 17134
rect 23940 17070 23992 17076
rect 23848 16788 23900 16794
rect 23848 16730 23900 16736
rect 23756 16516 23808 16522
rect 23756 16458 23808 16464
rect 23664 16448 23716 16454
rect 23664 16390 23716 16396
rect 23572 15428 23624 15434
rect 23572 15370 23624 15376
rect 23584 14958 23612 15370
rect 23768 15026 23796 16458
rect 23952 16046 23980 17070
rect 24110 16892 24418 16912
rect 24110 16890 24116 16892
rect 24172 16890 24196 16892
rect 24252 16890 24276 16892
rect 24332 16890 24356 16892
rect 24412 16890 24418 16892
rect 24172 16838 24174 16890
rect 24354 16838 24356 16890
rect 24110 16836 24116 16838
rect 24172 16836 24196 16838
rect 24252 16836 24276 16838
rect 24332 16836 24356 16838
rect 24412 16836 24418 16838
rect 24110 16816 24418 16836
rect 24584 16516 24636 16522
rect 24584 16458 24636 16464
rect 24596 16250 24624 16458
rect 24584 16244 24636 16250
rect 24584 16186 24636 16192
rect 24688 16130 24716 19246
rect 25056 16794 25084 21626
rect 28092 21146 28120 26930
rect 28354 26616 28410 26625
rect 28354 26551 28356 26560
rect 28408 26551 28410 26560
rect 28356 26522 28408 26528
rect 28356 25288 28408 25294
rect 28354 25256 28356 25265
rect 28408 25256 28410 25265
rect 28354 25191 28410 25200
rect 28172 25152 28224 25158
rect 28172 25094 28224 25100
rect 28080 21140 28132 21146
rect 28080 21082 28132 21088
rect 25412 17536 25464 17542
rect 25412 17478 25464 17484
rect 25424 17338 25452 17478
rect 25412 17332 25464 17338
rect 25412 17274 25464 17280
rect 25044 16788 25096 16794
rect 25044 16730 25096 16736
rect 25056 16590 25084 16730
rect 25044 16584 25096 16590
rect 25044 16526 25096 16532
rect 24596 16102 24716 16130
rect 26424 16108 26476 16114
rect 23940 16040 23992 16046
rect 23940 15982 23992 15988
rect 23848 15700 23900 15706
rect 23848 15642 23900 15648
rect 23860 15201 23888 15642
rect 23952 15570 23980 15982
rect 24110 15804 24418 15824
rect 24110 15802 24116 15804
rect 24172 15802 24196 15804
rect 24252 15802 24276 15804
rect 24332 15802 24356 15804
rect 24412 15802 24418 15804
rect 24172 15750 24174 15802
rect 24354 15750 24356 15802
rect 24110 15748 24116 15750
rect 24172 15748 24196 15750
rect 24252 15748 24276 15750
rect 24332 15748 24356 15750
rect 24412 15748 24418 15750
rect 24110 15728 24418 15748
rect 23940 15564 23992 15570
rect 23940 15506 23992 15512
rect 23940 15360 23992 15366
rect 23940 15302 23992 15308
rect 23846 15192 23902 15201
rect 23846 15127 23902 15136
rect 23952 15094 23980 15302
rect 23940 15088 23992 15094
rect 23940 15030 23992 15036
rect 23756 15020 23808 15026
rect 23756 14962 23808 14968
rect 23572 14952 23624 14958
rect 23478 14920 23534 14929
rect 23572 14894 23624 14900
rect 23478 14855 23534 14864
rect 23492 14618 23520 14855
rect 24032 14816 24084 14822
rect 24032 14758 24084 14764
rect 23480 14612 23532 14618
rect 23480 14554 23532 14560
rect 23388 14272 23440 14278
rect 23388 14214 23440 14220
rect 23400 14006 23428 14214
rect 23388 14000 23440 14006
rect 23388 13942 23440 13948
rect 23492 13954 23520 14554
rect 24044 14550 24072 14758
rect 24110 14716 24418 14736
rect 24110 14714 24116 14716
rect 24172 14714 24196 14716
rect 24252 14714 24276 14716
rect 24332 14714 24356 14716
rect 24412 14714 24418 14716
rect 24172 14662 24174 14714
rect 24354 14662 24356 14714
rect 24110 14660 24116 14662
rect 24172 14660 24196 14662
rect 24252 14660 24276 14662
rect 24332 14660 24356 14662
rect 24412 14660 24418 14662
rect 24110 14640 24418 14660
rect 24032 14544 24084 14550
rect 24032 14486 24084 14492
rect 23848 14408 23900 14414
rect 23848 14350 23900 14356
rect 23940 14408 23992 14414
rect 23940 14350 23992 14356
rect 23492 13938 23612 13954
rect 23492 13932 23624 13938
rect 23492 13926 23572 13932
rect 23572 13874 23624 13880
rect 23388 13796 23440 13802
rect 23388 13738 23440 13744
rect 23400 13394 23428 13738
rect 23664 13728 23716 13734
rect 23664 13670 23716 13676
rect 23388 13388 23440 13394
rect 23388 13330 23440 13336
rect 23676 13326 23704 13670
rect 23860 13530 23888 14350
rect 23952 13870 23980 14350
rect 23940 13864 23992 13870
rect 23940 13806 23992 13812
rect 23848 13524 23900 13530
rect 23848 13466 23900 13472
rect 23952 13326 23980 13806
rect 23296 13320 23348 13326
rect 23296 13262 23348 13268
rect 23664 13320 23716 13326
rect 23664 13262 23716 13268
rect 23940 13320 23992 13326
rect 23940 13262 23992 13268
rect 24044 12986 24072 14486
rect 24492 14272 24544 14278
rect 24492 14214 24544 14220
rect 24504 13938 24532 14214
rect 24492 13932 24544 13938
rect 24492 13874 24544 13880
rect 24110 13628 24418 13648
rect 24110 13626 24116 13628
rect 24172 13626 24196 13628
rect 24252 13626 24276 13628
rect 24332 13626 24356 13628
rect 24412 13626 24418 13628
rect 24172 13574 24174 13626
rect 24354 13574 24356 13626
rect 24110 13572 24116 13574
rect 24172 13572 24196 13574
rect 24252 13572 24276 13574
rect 24332 13572 24356 13574
rect 24412 13572 24418 13574
rect 24110 13552 24418 13572
rect 24032 12980 24084 12986
rect 24032 12922 24084 12928
rect 23020 12844 23072 12850
rect 23020 12786 23072 12792
rect 22848 12406 22968 12434
rect 22836 8968 22888 8974
rect 22836 8910 22888 8916
rect 22848 8566 22876 8910
rect 22652 8560 22704 8566
rect 22652 8502 22704 8508
rect 22836 8560 22888 8566
rect 22836 8502 22888 8508
rect 22284 8084 22336 8090
rect 22284 8026 22336 8032
rect 22296 7342 22324 8026
rect 22652 7744 22704 7750
rect 22652 7686 22704 7692
rect 22664 7478 22692 7686
rect 22652 7472 22704 7478
rect 22652 7414 22704 7420
rect 22848 7342 22876 8502
rect 22284 7336 22336 7342
rect 22284 7278 22336 7284
rect 22836 7336 22888 7342
rect 22836 7278 22888 7284
rect 22848 7206 22876 7278
rect 22836 7200 22888 7206
rect 22836 7142 22888 7148
rect 22940 7018 22968 12406
rect 23032 11898 23060 12786
rect 23480 12640 23532 12646
rect 23480 12582 23532 12588
rect 23756 12640 23808 12646
rect 23756 12582 23808 12588
rect 23020 11892 23072 11898
rect 23020 11834 23072 11840
rect 23492 11762 23520 12582
rect 23768 12238 23796 12582
rect 24110 12540 24418 12560
rect 24110 12538 24116 12540
rect 24172 12538 24196 12540
rect 24252 12538 24276 12540
rect 24332 12538 24356 12540
rect 24412 12538 24418 12540
rect 24172 12486 24174 12538
rect 24354 12486 24356 12538
rect 24110 12484 24116 12486
rect 24172 12484 24196 12486
rect 24252 12484 24276 12486
rect 24332 12484 24356 12486
rect 24412 12484 24418 12486
rect 24110 12464 24418 12484
rect 23940 12436 23992 12442
rect 23940 12378 23992 12384
rect 23572 12232 23624 12238
rect 23572 12174 23624 12180
rect 23756 12232 23808 12238
rect 23756 12174 23808 12180
rect 23584 12102 23612 12174
rect 23572 12096 23624 12102
rect 23572 12038 23624 12044
rect 23480 11756 23532 11762
rect 23480 11698 23532 11704
rect 23492 10674 23520 11698
rect 23572 11552 23624 11558
rect 23572 11494 23624 11500
rect 23584 11218 23612 11494
rect 23572 11212 23624 11218
rect 23572 11154 23624 11160
rect 23480 10668 23532 10674
rect 23480 10610 23532 10616
rect 23020 10464 23072 10470
rect 23020 10406 23072 10412
rect 23032 9994 23060 10406
rect 23492 10062 23520 10610
rect 23768 10062 23796 12174
rect 23848 12096 23900 12102
rect 23848 12038 23900 12044
rect 23860 10742 23888 12038
rect 23848 10736 23900 10742
rect 23848 10678 23900 10684
rect 23480 10056 23532 10062
rect 23480 9998 23532 10004
rect 23756 10056 23808 10062
rect 23756 9998 23808 10004
rect 23020 9988 23072 9994
rect 23020 9930 23072 9936
rect 23492 9738 23520 9998
rect 23400 9710 23520 9738
rect 23400 9586 23428 9710
rect 23388 9580 23440 9586
rect 23388 9522 23440 9528
rect 23664 9376 23716 9382
rect 23664 9318 23716 9324
rect 23480 8424 23532 8430
rect 23480 8366 23532 8372
rect 23492 7886 23520 8366
rect 23676 7886 23704 9318
rect 23756 8492 23808 8498
rect 23756 8434 23808 8440
rect 23768 8090 23796 8434
rect 23756 8084 23808 8090
rect 23756 8026 23808 8032
rect 23952 7970 23980 12378
rect 24032 12232 24084 12238
rect 24032 12174 24084 12180
rect 24044 11286 24072 12174
rect 24504 11898 24532 13874
rect 24596 12918 24624 16102
rect 26424 16050 26476 16056
rect 25136 15496 25188 15502
rect 25136 15438 25188 15444
rect 25148 15162 25176 15438
rect 25136 15156 25188 15162
rect 25136 15098 25188 15104
rect 24860 15088 24912 15094
rect 24858 15056 24860 15065
rect 24912 15056 24914 15065
rect 24858 14991 24914 15000
rect 26056 14612 26108 14618
rect 26056 14554 26108 14560
rect 25872 14340 25924 14346
rect 25872 14282 25924 14288
rect 25884 14074 25912 14282
rect 26068 14074 26096 14554
rect 26436 14074 26464 16050
rect 28184 15706 28212 25094
rect 28356 23520 28408 23526
rect 28356 23462 28408 23468
rect 28368 23225 28396 23462
rect 28354 23216 28410 23225
rect 28354 23151 28410 23160
rect 28356 17196 28408 17202
rect 28356 17138 28408 17144
rect 28368 17105 28396 17138
rect 28354 17096 28410 17105
rect 28354 17031 28410 17040
rect 28356 16652 28408 16658
rect 28356 16594 28408 16600
rect 28368 16425 28396 16594
rect 28354 16416 28410 16425
rect 28354 16351 28410 16360
rect 28172 15700 28224 15706
rect 28172 15642 28224 15648
rect 28356 15496 28408 15502
rect 28356 15438 28408 15444
rect 28368 15065 28396 15438
rect 28354 15056 28410 15065
rect 28354 14991 28410 15000
rect 28080 14272 28132 14278
rect 28080 14214 28132 14220
rect 25872 14068 25924 14074
rect 25872 14010 25924 14016
rect 26056 14068 26108 14074
rect 26056 14010 26108 14016
rect 26424 14068 26476 14074
rect 26424 14010 26476 14016
rect 24952 13932 25004 13938
rect 24952 13874 25004 13880
rect 24676 13864 24728 13870
rect 24676 13806 24728 13812
rect 24688 13258 24716 13806
rect 24964 13530 24992 13874
rect 25044 13864 25096 13870
rect 25044 13806 25096 13812
rect 24952 13524 25004 13530
rect 24952 13466 25004 13472
rect 24858 13424 24914 13433
rect 24858 13359 24914 13368
rect 24952 13388 25004 13394
rect 24768 13320 24820 13326
rect 24768 13262 24820 13268
rect 24676 13252 24728 13258
rect 24676 13194 24728 13200
rect 24584 12912 24636 12918
rect 24584 12854 24636 12860
rect 24584 12640 24636 12646
rect 24584 12582 24636 12588
rect 24596 12238 24624 12582
rect 24688 12306 24716 13194
rect 24676 12300 24728 12306
rect 24676 12242 24728 12248
rect 24780 12238 24808 13262
rect 24872 13190 24900 13359
rect 24952 13330 25004 13336
rect 24860 13184 24912 13190
rect 24860 13126 24912 13132
rect 24964 12782 24992 13330
rect 24860 12776 24912 12782
rect 24860 12718 24912 12724
rect 24952 12776 25004 12782
rect 24952 12718 25004 12724
rect 24584 12232 24636 12238
rect 24584 12174 24636 12180
rect 24768 12232 24820 12238
rect 24768 12174 24820 12180
rect 24492 11892 24544 11898
rect 24492 11834 24544 11840
rect 24780 11830 24808 12174
rect 24872 11898 24900 12718
rect 25056 12374 25084 13806
rect 25412 13728 25464 13734
rect 25412 13670 25464 13676
rect 25320 13184 25372 13190
rect 25320 13126 25372 13132
rect 25044 12368 25096 12374
rect 25044 12310 25096 12316
rect 24860 11892 24912 11898
rect 24860 11834 24912 11840
rect 25332 11830 25360 13126
rect 25424 12850 25452 13670
rect 25596 13252 25648 13258
rect 25596 13194 25648 13200
rect 25608 12986 25636 13194
rect 25872 13184 25924 13190
rect 25872 13126 25924 13132
rect 25596 12980 25648 12986
rect 25596 12922 25648 12928
rect 25412 12844 25464 12850
rect 25412 12786 25464 12792
rect 25688 12640 25740 12646
rect 25688 12582 25740 12588
rect 25700 12170 25728 12582
rect 25688 12164 25740 12170
rect 25688 12106 25740 12112
rect 25780 12096 25832 12102
rect 25780 12038 25832 12044
rect 24768 11824 24820 11830
rect 24768 11766 24820 11772
rect 25320 11824 25372 11830
rect 25320 11766 25372 11772
rect 25136 11756 25188 11762
rect 25136 11698 25188 11704
rect 25044 11552 25096 11558
rect 25044 11494 25096 11500
rect 24110 11452 24418 11472
rect 24110 11450 24116 11452
rect 24172 11450 24196 11452
rect 24252 11450 24276 11452
rect 24332 11450 24356 11452
rect 24412 11450 24418 11452
rect 24172 11398 24174 11450
rect 24354 11398 24356 11450
rect 24110 11396 24116 11398
rect 24172 11396 24196 11398
rect 24252 11396 24276 11398
rect 24332 11396 24356 11398
rect 24412 11396 24418 11398
rect 24110 11376 24418 11396
rect 24032 11280 24084 11286
rect 24032 11222 24084 11228
rect 25056 11218 25084 11494
rect 25044 11212 25096 11218
rect 25044 11154 25096 11160
rect 25148 11150 25176 11698
rect 25504 11688 25556 11694
rect 25504 11630 25556 11636
rect 24952 11144 25004 11150
rect 24952 11086 25004 11092
rect 25136 11144 25188 11150
rect 25136 11086 25188 11092
rect 24676 10464 24728 10470
rect 24676 10406 24728 10412
rect 24110 10364 24418 10384
rect 24110 10362 24116 10364
rect 24172 10362 24196 10364
rect 24252 10362 24276 10364
rect 24332 10362 24356 10364
rect 24412 10362 24418 10364
rect 24172 10310 24174 10362
rect 24354 10310 24356 10362
rect 24110 10308 24116 10310
rect 24172 10308 24196 10310
rect 24252 10308 24276 10310
rect 24332 10308 24356 10310
rect 24412 10308 24418 10310
rect 24110 10288 24418 10308
rect 24492 9988 24544 9994
rect 24492 9930 24544 9936
rect 24032 9920 24084 9926
rect 24032 9862 24084 9868
rect 24044 9722 24072 9862
rect 24032 9716 24084 9722
rect 24032 9658 24084 9664
rect 24032 9444 24084 9450
rect 24032 9386 24084 9392
rect 23768 7942 23980 7970
rect 23480 7880 23532 7886
rect 23664 7880 23716 7886
rect 23532 7828 23612 7834
rect 23480 7822 23612 7828
rect 23664 7822 23716 7828
rect 23492 7806 23612 7822
rect 23584 7274 23612 7806
rect 23572 7268 23624 7274
rect 23572 7210 23624 7216
rect 23112 7200 23164 7206
rect 23112 7142 23164 7148
rect 22848 6990 22968 7018
rect 22100 6860 22152 6866
rect 22100 6802 22152 6808
rect 21640 6724 21692 6730
rect 21640 6666 21692 6672
rect 22008 6724 22060 6730
rect 22008 6666 22060 6672
rect 21652 5302 21680 6666
rect 22020 6322 22048 6666
rect 22008 6316 22060 6322
rect 22008 6258 22060 6264
rect 21824 6112 21876 6118
rect 22020 6100 22048 6258
rect 21876 6072 22048 6100
rect 22192 6112 22244 6118
rect 21824 6054 21876 6060
rect 22192 6054 22244 6060
rect 21836 5846 21864 6054
rect 22204 5914 22232 6054
rect 22192 5908 22244 5914
rect 22192 5850 22244 5856
rect 21824 5840 21876 5846
rect 21824 5782 21876 5788
rect 22100 5704 22152 5710
rect 22020 5652 22100 5658
rect 22020 5646 22152 5652
rect 22652 5704 22704 5710
rect 22652 5646 22704 5652
rect 22020 5630 22140 5646
rect 22020 5370 22048 5630
rect 22560 5568 22612 5574
rect 22560 5510 22612 5516
rect 22008 5364 22060 5370
rect 22008 5306 22060 5312
rect 21640 5296 21692 5302
rect 21640 5238 21692 5244
rect 21916 5228 21968 5234
rect 21916 5170 21968 5176
rect 21548 5160 21600 5166
rect 21548 5102 21600 5108
rect 21560 4622 21588 5102
rect 21928 4690 21956 5170
rect 21916 4684 21968 4690
rect 21916 4626 21968 4632
rect 21548 4616 21600 4622
rect 21548 4558 21600 4564
rect 21560 4282 21588 4558
rect 21824 4548 21876 4554
rect 21824 4490 21876 4496
rect 21548 4276 21600 4282
rect 21548 4218 21600 4224
rect 21836 4026 21864 4490
rect 21928 4214 21956 4626
rect 22020 4554 22048 5306
rect 22572 4622 22600 5510
rect 22664 5302 22692 5646
rect 22652 5296 22704 5302
rect 22652 5238 22704 5244
rect 22560 4616 22612 4622
rect 22560 4558 22612 4564
rect 22744 4616 22796 4622
rect 22744 4558 22796 4564
rect 22008 4548 22060 4554
rect 22008 4490 22060 4496
rect 21916 4208 21968 4214
rect 21916 4150 21968 4156
rect 22756 4078 22784 4558
rect 21916 4072 21968 4078
rect 21836 4020 21916 4026
rect 21836 4014 21968 4020
rect 22744 4072 22796 4078
rect 22744 4014 22796 4020
rect 21836 3998 21956 4014
rect 21928 3738 21956 3998
rect 21916 3732 21968 3738
rect 21916 3674 21968 3680
rect 21456 3528 21508 3534
rect 21456 3470 21508 3476
rect 22848 3466 22876 6990
rect 22928 6724 22980 6730
rect 22928 6666 22980 6672
rect 22940 6390 22968 6666
rect 22928 6384 22980 6390
rect 22928 6326 22980 6332
rect 23124 6322 23152 7142
rect 23584 6730 23612 7210
rect 23572 6724 23624 6730
rect 23572 6666 23624 6672
rect 23388 6656 23440 6662
rect 23388 6598 23440 6604
rect 23400 6322 23428 6598
rect 23112 6316 23164 6322
rect 23112 6258 23164 6264
rect 23388 6316 23440 6322
rect 23388 6258 23440 6264
rect 23020 6248 23072 6254
rect 23020 6190 23072 6196
rect 23032 5574 23060 6190
rect 23020 5568 23072 5574
rect 23020 5510 23072 5516
rect 23020 5228 23072 5234
rect 23020 5170 23072 5176
rect 23032 4690 23060 5170
rect 23584 5166 23612 6666
rect 23768 5846 23796 7942
rect 23940 7880 23992 7886
rect 23940 7822 23992 7828
rect 23952 7002 23980 7822
rect 24044 7546 24072 9386
rect 24110 9276 24418 9296
rect 24110 9274 24116 9276
rect 24172 9274 24196 9276
rect 24252 9274 24276 9276
rect 24332 9274 24356 9276
rect 24412 9274 24418 9276
rect 24172 9222 24174 9274
rect 24354 9222 24356 9274
rect 24110 9220 24116 9222
rect 24172 9220 24196 9222
rect 24252 9220 24276 9222
rect 24332 9220 24356 9222
rect 24412 9220 24418 9222
rect 24110 9200 24418 9220
rect 24110 8188 24418 8208
rect 24110 8186 24116 8188
rect 24172 8186 24196 8188
rect 24252 8186 24276 8188
rect 24332 8186 24356 8188
rect 24412 8186 24418 8188
rect 24172 8134 24174 8186
rect 24354 8134 24356 8186
rect 24110 8132 24116 8134
rect 24172 8132 24196 8134
rect 24252 8132 24276 8134
rect 24332 8132 24356 8134
rect 24412 8132 24418 8134
rect 24110 8112 24418 8132
rect 24032 7540 24084 7546
rect 24032 7482 24084 7488
rect 24504 7478 24532 9930
rect 24688 9722 24716 10406
rect 24676 9716 24728 9722
rect 24676 9658 24728 9664
rect 24964 9654 24992 11086
rect 25148 10538 25176 11086
rect 25516 10606 25544 11630
rect 25792 11150 25820 12038
rect 25780 11144 25832 11150
rect 25780 11086 25832 11092
rect 25504 10600 25556 10606
rect 25504 10542 25556 10548
rect 25688 10600 25740 10606
rect 25688 10542 25740 10548
rect 25136 10532 25188 10538
rect 25136 10474 25188 10480
rect 25516 10130 25544 10542
rect 25700 10266 25728 10542
rect 25688 10260 25740 10266
rect 25688 10202 25740 10208
rect 25504 10124 25556 10130
rect 25504 10066 25556 10072
rect 25136 9920 25188 9926
rect 25136 9862 25188 9868
rect 25148 9722 25176 9862
rect 25136 9716 25188 9722
rect 25136 9658 25188 9664
rect 25700 9654 25728 10202
rect 25792 10062 25820 11086
rect 25780 10056 25832 10062
rect 25780 9998 25832 10004
rect 24952 9648 25004 9654
rect 24952 9590 25004 9596
rect 25688 9648 25740 9654
rect 25688 9590 25740 9596
rect 24860 9512 24912 9518
rect 24860 9454 24912 9460
rect 24872 9042 24900 9454
rect 24964 9450 24992 9590
rect 24952 9444 25004 9450
rect 24952 9386 25004 9392
rect 24860 9036 24912 9042
rect 24860 8978 24912 8984
rect 24492 7472 24544 7478
rect 24492 7414 24544 7420
rect 24872 7410 24900 8978
rect 24964 7478 24992 9386
rect 25884 8922 25912 13126
rect 26056 12844 26108 12850
rect 26056 12786 26108 12792
rect 26068 12442 26096 12786
rect 26056 12436 26108 12442
rect 26056 12378 26108 12384
rect 25964 12096 26016 12102
rect 25964 12038 26016 12044
rect 25976 11898 26004 12038
rect 25964 11892 26016 11898
rect 25964 11834 26016 11840
rect 26056 11688 26108 11694
rect 26056 11630 26108 11636
rect 26068 11098 26096 11630
rect 26516 11348 26568 11354
rect 26516 11290 26568 11296
rect 26332 11144 26384 11150
rect 26068 11092 26332 11098
rect 26068 11086 26384 11092
rect 26068 11070 26372 11086
rect 26424 11076 26476 11082
rect 26068 9654 26096 11070
rect 26424 11018 26476 11024
rect 26436 10810 26464 11018
rect 26424 10804 26476 10810
rect 26424 10746 26476 10752
rect 26528 10674 26556 11290
rect 28092 10674 28120 14214
rect 28264 13932 28316 13938
rect 28264 13874 28316 13880
rect 28276 13705 28304 13874
rect 28262 13696 28318 13705
rect 28262 13631 28318 13640
rect 28356 12640 28408 12646
rect 28356 12582 28408 12588
rect 28368 12345 28396 12582
rect 28354 12336 28410 12345
rect 28354 12271 28410 12280
rect 28264 11756 28316 11762
rect 28264 11698 28316 11704
rect 28276 11665 28304 11698
rect 28262 11656 28318 11665
rect 28262 11591 28318 11600
rect 26516 10668 26568 10674
rect 26516 10610 26568 10616
rect 28080 10668 28132 10674
rect 28080 10610 28132 10616
rect 26148 10464 26200 10470
rect 26148 10406 26200 10412
rect 28264 10464 28316 10470
rect 28264 10406 28316 10412
rect 26160 9722 26188 10406
rect 28276 10305 28304 10406
rect 28262 10296 28318 10305
rect 28262 10231 28318 10240
rect 27436 10056 27488 10062
rect 27436 9998 27488 10004
rect 27448 9722 27476 9998
rect 26148 9716 26200 9722
rect 26148 9658 26200 9664
rect 27436 9716 27488 9722
rect 27436 9658 27488 9664
rect 26056 9648 26108 9654
rect 26056 9590 26108 9596
rect 28356 8968 28408 8974
rect 25792 8894 25912 8922
rect 28354 8936 28356 8945
rect 28408 8936 28410 8945
rect 25136 8832 25188 8838
rect 25136 8774 25188 8780
rect 25228 8832 25280 8838
rect 25228 8774 25280 8780
rect 25148 8090 25176 8774
rect 25240 8634 25268 8774
rect 25228 8628 25280 8634
rect 25228 8570 25280 8576
rect 25136 8084 25188 8090
rect 25136 8026 25188 8032
rect 25240 7546 25268 8570
rect 25412 7880 25464 7886
rect 25412 7822 25464 7828
rect 25228 7540 25280 7546
rect 25228 7482 25280 7488
rect 24952 7472 25004 7478
rect 24952 7414 25004 7420
rect 24860 7404 24912 7410
rect 24860 7346 24912 7352
rect 24110 7100 24418 7120
rect 24110 7098 24116 7100
rect 24172 7098 24196 7100
rect 24252 7098 24276 7100
rect 24332 7098 24356 7100
rect 24412 7098 24418 7100
rect 24172 7046 24174 7098
rect 24354 7046 24356 7098
rect 24110 7044 24116 7046
rect 24172 7044 24196 7046
rect 24252 7044 24276 7046
rect 24332 7044 24356 7046
rect 24412 7044 24418 7046
rect 24110 7024 24418 7044
rect 23940 6996 23992 7002
rect 23940 6938 23992 6944
rect 23952 6458 23980 6938
rect 24676 6724 24728 6730
rect 24676 6666 24728 6672
rect 23940 6452 23992 6458
rect 23940 6394 23992 6400
rect 24688 6322 24716 6666
rect 23848 6316 23900 6322
rect 23848 6258 23900 6264
rect 24676 6316 24728 6322
rect 24676 6258 24728 6264
rect 23860 5914 23888 6258
rect 24032 6112 24084 6118
rect 24032 6054 24084 6060
rect 23848 5908 23900 5914
rect 23848 5850 23900 5856
rect 23756 5840 23808 5846
rect 23756 5782 23808 5788
rect 23768 5710 23796 5782
rect 23756 5704 23808 5710
rect 23756 5646 23808 5652
rect 24044 5302 24072 6054
rect 24110 6012 24418 6032
rect 24110 6010 24116 6012
rect 24172 6010 24196 6012
rect 24252 6010 24276 6012
rect 24332 6010 24356 6012
rect 24412 6010 24418 6012
rect 24172 5958 24174 6010
rect 24354 5958 24356 6010
rect 24110 5956 24116 5958
rect 24172 5956 24196 5958
rect 24252 5956 24276 5958
rect 24332 5956 24356 5958
rect 24412 5956 24418 5958
rect 24110 5936 24418 5956
rect 24688 5778 24716 6258
rect 24872 6186 24900 7346
rect 24964 6934 24992 7414
rect 25320 7200 25372 7206
rect 25320 7142 25372 7148
rect 24952 6928 25004 6934
rect 24952 6870 25004 6876
rect 25136 6656 25188 6662
rect 25136 6598 25188 6604
rect 25148 6322 25176 6598
rect 25332 6390 25360 7142
rect 25424 6390 25452 7822
rect 25792 7750 25820 8894
rect 28354 8871 28410 8880
rect 25872 8832 25924 8838
rect 25872 8774 25924 8780
rect 25884 8566 25912 8774
rect 25872 8560 25924 8566
rect 25872 8502 25924 8508
rect 26148 8288 26200 8294
rect 26148 8230 26200 8236
rect 25872 7948 25924 7954
rect 25872 7890 25924 7896
rect 25780 7744 25832 7750
rect 25780 7686 25832 7692
rect 25884 7342 25912 7890
rect 26160 7886 26188 8230
rect 26148 7880 26200 7886
rect 26148 7822 26200 7828
rect 28356 7880 28408 7886
rect 28356 7822 28408 7828
rect 28368 7585 28396 7822
rect 28354 7576 28410 7585
rect 28354 7511 28410 7520
rect 25872 7336 25924 7342
rect 25872 7278 25924 7284
rect 25688 6724 25740 6730
rect 25688 6666 25740 6672
rect 25700 6458 25728 6666
rect 25688 6452 25740 6458
rect 25688 6394 25740 6400
rect 25320 6384 25372 6390
rect 25320 6326 25372 6332
rect 25412 6384 25464 6390
rect 25412 6326 25464 6332
rect 25136 6316 25188 6322
rect 25136 6258 25188 6264
rect 24860 6180 24912 6186
rect 24860 6122 24912 6128
rect 24676 5772 24728 5778
rect 24676 5714 24728 5720
rect 24032 5296 24084 5302
rect 24032 5238 24084 5244
rect 24872 5234 24900 6122
rect 25148 5710 25176 6258
rect 25136 5704 25188 5710
rect 25136 5646 25188 5652
rect 28356 5704 28408 5710
rect 28356 5646 28408 5652
rect 25228 5568 25280 5574
rect 28368 5545 28396 5646
rect 25228 5510 25280 5516
rect 28354 5536 28410 5545
rect 24860 5228 24912 5234
rect 24860 5170 24912 5176
rect 23572 5160 23624 5166
rect 23572 5102 23624 5108
rect 25240 5030 25268 5510
rect 28354 5471 28410 5480
rect 23112 5024 23164 5030
rect 23112 4966 23164 4972
rect 24492 5024 24544 5030
rect 24492 4966 24544 4972
rect 25228 5024 25280 5030
rect 25228 4966 25280 4972
rect 23124 4826 23152 4966
rect 24110 4924 24418 4944
rect 24110 4922 24116 4924
rect 24172 4922 24196 4924
rect 24252 4922 24276 4924
rect 24332 4922 24356 4924
rect 24412 4922 24418 4924
rect 24172 4870 24174 4922
rect 24354 4870 24356 4922
rect 24110 4868 24116 4870
rect 24172 4868 24196 4870
rect 24252 4868 24276 4870
rect 24332 4868 24356 4870
rect 24412 4868 24418 4870
rect 24110 4848 24418 4868
rect 23112 4820 23164 4826
rect 23112 4762 23164 4768
rect 23940 4752 23992 4758
rect 23940 4694 23992 4700
rect 23020 4684 23072 4690
rect 23020 4626 23072 4632
rect 23952 4146 23980 4694
rect 23940 4140 23992 4146
rect 23940 4082 23992 4088
rect 24504 4078 24532 4966
rect 24492 4072 24544 4078
rect 24492 4014 24544 4020
rect 24110 3836 24418 3856
rect 24110 3834 24116 3836
rect 24172 3834 24196 3836
rect 24252 3834 24276 3836
rect 24332 3834 24356 3836
rect 24412 3834 24418 3836
rect 24172 3782 24174 3834
rect 24354 3782 24356 3834
rect 24110 3780 24116 3782
rect 24172 3780 24196 3782
rect 24252 3780 24276 3782
rect 24332 3780 24356 3782
rect 24412 3780 24418 3782
rect 24110 3760 24418 3780
rect 24504 3534 24532 4014
rect 24492 3528 24544 3534
rect 24492 3470 24544 3476
rect 22836 3460 22888 3466
rect 22836 3402 22888 3408
rect 22284 3392 22336 3398
rect 22284 3334 22336 3340
rect 20720 2644 20772 2650
rect 20720 2586 20772 2592
rect 20444 2576 20496 2582
rect 20444 2518 20496 2524
rect 18512 2508 18564 2514
rect 18512 2450 18564 2456
rect 20352 2508 20404 2514
rect 20352 2450 20404 2456
rect 22296 2446 22324 3334
rect 24110 2748 24418 2768
rect 24110 2746 24116 2748
rect 24172 2746 24196 2748
rect 24252 2746 24276 2748
rect 24332 2746 24356 2748
rect 24412 2746 24418 2748
rect 24172 2694 24174 2746
rect 24354 2694 24356 2746
rect 24110 2692 24116 2694
rect 24172 2692 24196 2694
rect 24252 2692 24276 2694
rect 24332 2692 24356 2694
rect 24412 2692 24418 2694
rect 24110 2672 24418 2692
rect 25240 2446 25268 4966
rect 28356 4616 28408 4622
rect 28356 4558 28408 4564
rect 28368 4185 28396 4558
rect 28354 4176 28410 4185
rect 28354 4111 28410 4120
rect 28080 3392 28132 3398
rect 28080 3334 28132 3340
rect 28092 3058 28120 3334
rect 28080 3052 28132 3058
rect 28080 2994 28132 3000
rect 28264 2848 28316 2854
rect 28264 2790 28316 2796
rect 20720 2440 20772 2446
rect 20640 2400 20720 2428
rect 15660 2372 15712 2378
rect 15660 2314 15712 2320
rect 16764 2372 16816 2378
rect 16764 2314 16816 2320
rect 16776 800 16804 2314
rect 18696 2304 18748 2310
rect 18696 2246 18748 2252
rect 18708 800 18736 2246
rect 19478 2204 19786 2224
rect 19478 2202 19484 2204
rect 19540 2202 19564 2204
rect 19620 2202 19644 2204
rect 19700 2202 19724 2204
rect 19780 2202 19786 2204
rect 19540 2150 19542 2202
rect 19722 2150 19724 2202
rect 19478 2148 19484 2150
rect 19540 2148 19564 2150
rect 19620 2148 19644 2150
rect 19700 2148 19724 2150
rect 19780 2148 19786 2150
rect 19478 2128 19786 2148
rect 20640 800 20668 2400
rect 20720 2382 20772 2388
rect 22284 2440 22336 2446
rect 22284 2382 22336 2388
rect 25228 2440 25280 2446
rect 25228 2382 25280 2388
rect 26424 2440 26476 2446
rect 26424 2382 26476 2388
rect 21916 2304 21968 2310
rect 21916 2246 21968 2252
rect 25136 2304 25188 2310
rect 25136 2246 25188 2252
rect 21928 800 21956 2246
rect 25148 800 25176 2246
rect 26436 800 26464 2382
rect 27712 2304 27764 2310
rect 27712 2246 27764 2252
rect 27724 800 27752 2246
rect 1674 776 1730 785
rect 1674 711 1730 720
rect 1950 0 2006 800
rect 3238 0 3294 800
rect 3882 0 3938 800
rect 5170 0 5226 800
rect 6458 0 6514 800
rect 7746 0 7802 800
rect 8390 0 8446 800
rect 9678 0 9734 800
rect 10966 0 11022 800
rect 12254 0 12310 800
rect 12898 0 12954 800
rect 14186 0 14242 800
rect 15474 0 15530 800
rect 16762 0 16818 800
rect 17406 0 17462 800
rect 18694 0 18750 800
rect 19982 0 20038 800
rect 20626 0 20682 800
rect 21914 0 21970 800
rect 23202 0 23258 800
rect 24490 0 24546 800
rect 25134 0 25190 800
rect 26422 0 26478 800
rect 27710 0 27766 800
rect 28276 785 28304 2790
rect 28262 776 28318 785
rect 28262 711 28318 720
rect 28998 0 29054 800
rect 29642 0 29698 800
<< via2 >>
rect 1674 27920 1730 27976
rect 5588 27770 5644 27772
rect 5668 27770 5724 27772
rect 5748 27770 5804 27772
rect 5828 27770 5884 27772
rect 5588 27718 5634 27770
rect 5634 27718 5644 27770
rect 5668 27718 5698 27770
rect 5698 27718 5710 27770
rect 5710 27718 5724 27770
rect 5748 27718 5762 27770
rect 5762 27718 5774 27770
rect 5774 27718 5804 27770
rect 5828 27718 5838 27770
rect 5838 27718 5884 27770
rect 5588 27716 5644 27718
rect 5668 27716 5724 27718
rect 5748 27716 5804 27718
rect 5828 27716 5884 27718
rect 1398 26560 1454 26616
rect 1398 25880 1454 25936
rect 1398 24520 1454 24576
rect 1398 23160 1454 23216
rect 1398 21120 1454 21176
rect 1398 19796 1400 19816
rect 1400 19796 1452 19816
rect 1452 19796 1454 19816
rect 1398 19760 1454 19796
rect 1398 18400 1454 18456
rect 1398 17060 1454 17096
rect 1398 17040 1400 17060
rect 1400 17040 1452 17060
rect 1452 17040 1454 17060
rect 5588 26682 5644 26684
rect 5668 26682 5724 26684
rect 5748 26682 5804 26684
rect 5828 26682 5884 26684
rect 5588 26630 5634 26682
rect 5634 26630 5644 26682
rect 5668 26630 5698 26682
rect 5698 26630 5710 26682
rect 5710 26630 5724 26682
rect 5748 26630 5762 26682
rect 5762 26630 5774 26682
rect 5774 26630 5804 26682
rect 5828 26630 5838 26682
rect 5838 26630 5884 26682
rect 5588 26628 5644 26630
rect 5668 26628 5724 26630
rect 5748 26628 5804 26630
rect 5828 26628 5884 26630
rect 5588 25594 5644 25596
rect 5668 25594 5724 25596
rect 5748 25594 5804 25596
rect 5828 25594 5884 25596
rect 5588 25542 5634 25594
rect 5634 25542 5644 25594
rect 5668 25542 5698 25594
rect 5698 25542 5710 25594
rect 5710 25542 5724 25594
rect 5748 25542 5762 25594
rect 5762 25542 5774 25594
rect 5774 25542 5804 25594
rect 5828 25542 5838 25594
rect 5838 25542 5884 25594
rect 5588 25540 5644 25542
rect 5668 25540 5724 25542
rect 5748 25540 5804 25542
rect 5828 25540 5884 25542
rect 14852 27770 14908 27772
rect 14932 27770 14988 27772
rect 15012 27770 15068 27772
rect 15092 27770 15148 27772
rect 14852 27718 14898 27770
rect 14898 27718 14908 27770
rect 14932 27718 14962 27770
rect 14962 27718 14974 27770
rect 14974 27718 14988 27770
rect 15012 27718 15026 27770
rect 15026 27718 15038 27770
rect 15038 27718 15068 27770
rect 15092 27718 15102 27770
rect 15102 27718 15148 27770
rect 14852 27716 14908 27718
rect 14932 27716 14988 27718
rect 15012 27716 15068 27718
rect 15092 27716 15148 27718
rect 24116 27770 24172 27772
rect 24196 27770 24252 27772
rect 24276 27770 24332 27772
rect 24356 27770 24412 27772
rect 24116 27718 24162 27770
rect 24162 27718 24172 27770
rect 24196 27718 24226 27770
rect 24226 27718 24238 27770
rect 24238 27718 24252 27770
rect 24276 27718 24290 27770
rect 24290 27718 24302 27770
rect 24302 27718 24332 27770
rect 24356 27718 24366 27770
rect 24366 27718 24412 27770
rect 24116 27716 24172 27718
rect 24196 27716 24252 27718
rect 24276 27716 24332 27718
rect 24356 27716 24412 27718
rect 27526 29280 27582 29336
rect 10220 27226 10276 27228
rect 10300 27226 10356 27228
rect 10380 27226 10436 27228
rect 10460 27226 10516 27228
rect 10220 27174 10266 27226
rect 10266 27174 10276 27226
rect 10300 27174 10330 27226
rect 10330 27174 10342 27226
rect 10342 27174 10356 27226
rect 10380 27174 10394 27226
rect 10394 27174 10406 27226
rect 10406 27174 10436 27226
rect 10460 27174 10470 27226
rect 10470 27174 10516 27226
rect 10220 27172 10276 27174
rect 10300 27172 10356 27174
rect 10380 27172 10436 27174
rect 10460 27172 10516 27174
rect 10220 26138 10276 26140
rect 10300 26138 10356 26140
rect 10380 26138 10436 26140
rect 10460 26138 10516 26140
rect 10220 26086 10266 26138
rect 10266 26086 10276 26138
rect 10300 26086 10330 26138
rect 10330 26086 10342 26138
rect 10342 26086 10356 26138
rect 10380 26086 10394 26138
rect 10394 26086 10406 26138
rect 10406 26086 10436 26138
rect 10460 26086 10470 26138
rect 10470 26086 10516 26138
rect 10220 26084 10276 26086
rect 10300 26084 10356 26086
rect 10380 26084 10436 26086
rect 10460 26084 10516 26086
rect 10220 25050 10276 25052
rect 10300 25050 10356 25052
rect 10380 25050 10436 25052
rect 10460 25050 10516 25052
rect 10220 24998 10266 25050
rect 10266 24998 10276 25050
rect 10300 24998 10330 25050
rect 10330 24998 10342 25050
rect 10342 24998 10356 25050
rect 10380 24998 10394 25050
rect 10394 24998 10406 25050
rect 10406 24998 10436 25050
rect 10460 24998 10470 25050
rect 10470 24998 10516 25050
rect 10220 24996 10276 24998
rect 10300 24996 10356 24998
rect 10380 24996 10436 24998
rect 10460 24996 10516 24998
rect 5588 24506 5644 24508
rect 5668 24506 5724 24508
rect 5748 24506 5804 24508
rect 5828 24506 5884 24508
rect 5588 24454 5634 24506
rect 5634 24454 5644 24506
rect 5668 24454 5698 24506
rect 5698 24454 5710 24506
rect 5710 24454 5724 24506
rect 5748 24454 5762 24506
rect 5762 24454 5774 24506
rect 5774 24454 5804 24506
rect 5828 24454 5838 24506
rect 5838 24454 5884 24506
rect 5588 24452 5644 24454
rect 5668 24452 5724 24454
rect 5748 24452 5804 24454
rect 5828 24452 5884 24454
rect 10220 23962 10276 23964
rect 10300 23962 10356 23964
rect 10380 23962 10436 23964
rect 10460 23962 10516 23964
rect 10220 23910 10266 23962
rect 10266 23910 10276 23962
rect 10300 23910 10330 23962
rect 10330 23910 10342 23962
rect 10342 23910 10356 23962
rect 10380 23910 10394 23962
rect 10394 23910 10406 23962
rect 10406 23910 10436 23962
rect 10460 23910 10470 23962
rect 10470 23910 10516 23962
rect 10220 23908 10276 23910
rect 10300 23908 10356 23910
rect 10380 23908 10436 23910
rect 10460 23908 10516 23910
rect 5588 23418 5644 23420
rect 5668 23418 5724 23420
rect 5748 23418 5804 23420
rect 5828 23418 5884 23420
rect 5588 23366 5634 23418
rect 5634 23366 5644 23418
rect 5668 23366 5698 23418
rect 5698 23366 5710 23418
rect 5710 23366 5724 23418
rect 5748 23366 5762 23418
rect 5762 23366 5774 23418
rect 5774 23366 5804 23418
rect 5828 23366 5838 23418
rect 5838 23366 5884 23418
rect 5588 23364 5644 23366
rect 5668 23364 5724 23366
rect 5748 23364 5804 23366
rect 5828 23364 5884 23366
rect 10220 22874 10276 22876
rect 10300 22874 10356 22876
rect 10380 22874 10436 22876
rect 10460 22874 10516 22876
rect 10220 22822 10266 22874
rect 10266 22822 10276 22874
rect 10300 22822 10330 22874
rect 10330 22822 10342 22874
rect 10342 22822 10356 22874
rect 10380 22822 10394 22874
rect 10394 22822 10406 22874
rect 10406 22822 10436 22874
rect 10460 22822 10470 22874
rect 10470 22822 10516 22874
rect 10220 22820 10276 22822
rect 10300 22820 10356 22822
rect 10380 22820 10436 22822
rect 10460 22820 10516 22822
rect 5588 22330 5644 22332
rect 5668 22330 5724 22332
rect 5748 22330 5804 22332
rect 5828 22330 5884 22332
rect 5588 22278 5634 22330
rect 5634 22278 5644 22330
rect 5668 22278 5698 22330
rect 5698 22278 5710 22330
rect 5710 22278 5724 22330
rect 5748 22278 5762 22330
rect 5762 22278 5774 22330
rect 5774 22278 5804 22330
rect 5828 22278 5838 22330
rect 5838 22278 5884 22330
rect 5588 22276 5644 22278
rect 5668 22276 5724 22278
rect 5748 22276 5804 22278
rect 5828 22276 5884 22278
rect 5588 21242 5644 21244
rect 5668 21242 5724 21244
rect 5748 21242 5804 21244
rect 5828 21242 5884 21244
rect 5588 21190 5634 21242
rect 5634 21190 5644 21242
rect 5668 21190 5698 21242
rect 5698 21190 5710 21242
rect 5710 21190 5724 21242
rect 5748 21190 5762 21242
rect 5762 21190 5774 21242
rect 5774 21190 5804 21242
rect 5828 21190 5838 21242
rect 5838 21190 5884 21242
rect 5588 21188 5644 21190
rect 5668 21188 5724 21190
rect 5748 21188 5804 21190
rect 5828 21188 5884 21190
rect 5588 20154 5644 20156
rect 5668 20154 5724 20156
rect 5748 20154 5804 20156
rect 5828 20154 5884 20156
rect 5588 20102 5634 20154
rect 5634 20102 5644 20154
rect 5668 20102 5698 20154
rect 5698 20102 5710 20154
rect 5710 20102 5724 20154
rect 5748 20102 5762 20154
rect 5762 20102 5774 20154
rect 5774 20102 5804 20154
rect 5828 20102 5838 20154
rect 5838 20102 5884 20154
rect 5588 20100 5644 20102
rect 5668 20100 5724 20102
rect 5748 20100 5804 20102
rect 5828 20100 5884 20102
rect 10220 21786 10276 21788
rect 10300 21786 10356 21788
rect 10380 21786 10436 21788
rect 10460 21786 10516 21788
rect 10220 21734 10266 21786
rect 10266 21734 10276 21786
rect 10300 21734 10330 21786
rect 10330 21734 10342 21786
rect 10342 21734 10356 21786
rect 10380 21734 10394 21786
rect 10394 21734 10406 21786
rect 10406 21734 10436 21786
rect 10460 21734 10470 21786
rect 10470 21734 10516 21786
rect 10220 21732 10276 21734
rect 10300 21732 10356 21734
rect 10380 21732 10436 21734
rect 10460 21732 10516 21734
rect 10220 20698 10276 20700
rect 10300 20698 10356 20700
rect 10380 20698 10436 20700
rect 10460 20698 10516 20700
rect 10220 20646 10266 20698
rect 10266 20646 10276 20698
rect 10300 20646 10330 20698
rect 10330 20646 10342 20698
rect 10342 20646 10356 20698
rect 10380 20646 10394 20698
rect 10394 20646 10406 20698
rect 10406 20646 10436 20698
rect 10460 20646 10470 20698
rect 10470 20646 10516 20698
rect 10220 20644 10276 20646
rect 10300 20644 10356 20646
rect 10380 20644 10436 20646
rect 10460 20644 10516 20646
rect 5588 19066 5644 19068
rect 5668 19066 5724 19068
rect 5748 19066 5804 19068
rect 5828 19066 5884 19068
rect 5588 19014 5634 19066
rect 5634 19014 5644 19066
rect 5668 19014 5698 19066
rect 5698 19014 5710 19066
rect 5710 19014 5724 19066
rect 5748 19014 5762 19066
rect 5762 19014 5774 19066
rect 5774 19014 5804 19066
rect 5828 19014 5838 19066
rect 5838 19014 5884 19066
rect 5588 19012 5644 19014
rect 5668 19012 5724 19014
rect 5748 19012 5804 19014
rect 5828 19012 5884 19014
rect 1766 17176 1822 17232
rect 5588 17978 5644 17980
rect 5668 17978 5724 17980
rect 5748 17978 5804 17980
rect 5828 17978 5884 17980
rect 5588 17926 5634 17978
rect 5634 17926 5644 17978
rect 5668 17926 5698 17978
rect 5698 17926 5710 17978
rect 5710 17926 5724 17978
rect 5748 17926 5762 17978
rect 5762 17926 5774 17978
rect 5774 17926 5804 17978
rect 5828 17926 5838 17978
rect 5838 17926 5884 17978
rect 5588 17924 5644 17926
rect 5668 17924 5724 17926
rect 5748 17924 5804 17926
rect 5828 17924 5884 17926
rect 5588 16890 5644 16892
rect 5668 16890 5724 16892
rect 5748 16890 5804 16892
rect 5828 16890 5884 16892
rect 5588 16838 5634 16890
rect 5634 16838 5644 16890
rect 5668 16838 5698 16890
rect 5698 16838 5710 16890
rect 5710 16838 5724 16890
rect 5748 16838 5762 16890
rect 5762 16838 5774 16890
rect 5774 16838 5804 16890
rect 5828 16838 5838 16890
rect 5838 16838 5884 16890
rect 5588 16836 5644 16838
rect 5668 16836 5724 16838
rect 5748 16836 5804 16838
rect 5828 16836 5884 16838
rect 1490 16396 1492 16416
rect 1492 16396 1544 16416
rect 1544 16396 1546 16416
rect 1490 16360 1546 16396
rect 1398 13640 1454 13696
rect 1398 10240 1454 10296
rect 1674 8900 1730 8936
rect 1674 8880 1676 8900
rect 1676 8880 1728 8900
rect 1728 8880 1730 8900
rect 5588 15802 5644 15804
rect 5668 15802 5724 15804
rect 5748 15802 5804 15804
rect 5828 15802 5884 15804
rect 5588 15750 5634 15802
rect 5634 15750 5644 15802
rect 5668 15750 5698 15802
rect 5698 15750 5710 15802
rect 5710 15750 5724 15802
rect 5748 15750 5762 15802
rect 5762 15750 5774 15802
rect 5774 15750 5804 15802
rect 5828 15750 5838 15802
rect 5838 15750 5884 15802
rect 5588 15748 5644 15750
rect 5668 15748 5724 15750
rect 5748 15748 5804 15750
rect 5828 15748 5884 15750
rect 5588 14714 5644 14716
rect 5668 14714 5724 14716
rect 5748 14714 5804 14716
rect 5828 14714 5884 14716
rect 5588 14662 5634 14714
rect 5634 14662 5644 14714
rect 5668 14662 5698 14714
rect 5698 14662 5710 14714
rect 5710 14662 5724 14714
rect 5748 14662 5762 14714
rect 5762 14662 5774 14714
rect 5774 14662 5804 14714
rect 5828 14662 5838 14714
rect 5838 14662 5884 14714
rect 5588 14660 5644 14662
rect 5668 14660 5724 14662
rect 5748 14660 5804 14662
rect 5828 14660 5884 14662
rect 5588 13626 5644 13628
rect 5668 13626 5724 13628
rect 5748 13626 5804 13628
rect 5828 13626 5884 13628
rect 5588 13574 5634 13626
rect 5634 13574 5644 13626
rect 5668 13574 5698 13626
rect 5698 13574 5710 13626
rect 5710 13574 5724 13626
rect 5748 13574 5762 13626
rect 5762 13574 5774 13626
rect 5774 13574 5804 13626
rect 5828 13574 5838 13626
rect 5838 13574 5884 13626
rect 5588 13572 5644 13574
rect 5668 13572 5724 13574
rect 5748 13572 5804 13574
rect 5828 13572 5884 13574
rect 5588 12538 5644 12540
rect 5668 12538 5724 12540
rect 5748 12538 5804 12540
rect 5828 12538 5884 12540
rect 5588 12486 5634 12538
rect 5634 12486 5644 12538
rect 5668 12486 5698 12538
rect 5698 12486 5710 12538
rect 5710 12486 5724 12538
rect 5748 12486 5762 12538
rect 5762 12486 5774 12538
rect 5774 12486 5804 12538
rect 5828 12486 5838 12538
rect 5838 12486 5884 12538
rect 5588 12484 5644 12486
rect 5668 12484 5724 12486
rect 5748 12484 5804 12486
rect 5828 12484 5884 12486
rect 5588 11450 5644 11452
rect 5668 11450 5724 11452
rect 5748 11450 5804 11452
rect 5828 11450 5884 11452
rect 5588 11398 5634 11450
rect 5634 11398 5644 11450
rect 5668 11398 5698 11450
rect 5698 11398 5710 11450
rect 5710 11398 5724 11450
rect 5748 11398 5762 11450
rect 5762 11398 5774 11450
rect 5774 11398 5804 11450
rect 5828 11398 5838 11450
rect 5838 11398 5884 11450
rect 5588 11396 5644 11398
rect 5668 11396 5724 11398
rect 5748 11396 5804 11398
rect 5828 11396 5884 11398
rect 5588 10362 5644 10364
rect 5668 10362 5724 10364
rect 5748 10362 5804 10364
rect 5828 10362 5884 10364
rect 5588 10310 5634 10362
rect 5634 10310 5644 10362
rect 5668 10310 5698 10362
rect 5698 10310 5710 10362
rect 5710 10310 5724 10362
rect 5748 10310 5762 10362
rect 5762 10310 5774 10362
rect 5774 10310 5804 10362
rect 5828 10310 5838 10362
rect 5838 10310 5884 10362
rect 5588 10308 5644 10310
rect 5668 10308 5724 10310
rect 5748 10308 5804 10310
rect 5828 10308 5884 10310
rect 10220 19610 10276 19612
rect 10300 19610 10356 19612
rect 10380 19610 10436 19612
rect 10460 19610 10516 19612
rect 10220 19558 10266 19610
rect 10266 19558 10276 19610
rect 10300 19558 10330 19610
rect 10330 19558 10342 19610
rect 10342 19558 10356 19610
rect 10380 19558 10394 19610
rect 10394 19558 10406 19610
rect 10406 19558 10436 19610
rect 10460 19558 10470 19610
rect 10470 19558 10516 19610
rect 10220 19556 10276 19558
rect 10300 19556 10356 19558
rect 10380 19556 10436 19558
rect 10460 19556 10516 19558
rect 10220 18522 10276 18524
rect 10300 18522 10356 18524
rect 10380 18522 10436 18524
rect 10460 18522 10516 18524
rect 10220 18470 10266 18522
rect 10266 18470 10276 18522
rect 10300 18470 10330 18522
rect 10330 18470 10342 18522
rect 10342 18470 10356 18522
rect 10380 18470 10394 18522
rect 10394 18470 10406 18522
rect 10406 18470 10436 18522
rect 10460 18470 10470 18522
rect 10470 18470 10516 18522
rect 10220 18468 10276 18470
rect 10300 18468 10356 18470
rect 10380 18468 10436 18470
rect 10460 18468 10516 18470
rect 10220 17434 10276 17436
rect 10300 17434 10356 17436
rect 10380 17434 10436 17436
rect 10460 17434 10516 17436
rect 10220 17382 10266 17434
rect 10266 17382 10276 17434
rect 10300 17382 10330 17434
rect 10330 17382 10342 17434
rect 10342 17382 10356 17434
rect 10380 17382 10394 17434
rect 10394 17382 10406 17434
rect 10406 17382 10436 17434
rect 10460 17382 10470 17434
rect 10470 17382 10516 17434
rect 10220 17380 10276 17382
rect 10300 17380 10356 17382
rect 10380 17380 10436 17382
rect 10460 17380 10516 17382
rect 14852 26682 14908 26684
rect 14932 26682 14988 26684
rect 15012 26682 15068 26684
rect 15092 26682 15148 26684
rect 14852 26630 14898 26682
rect 14898 26630 14908 26682
rect 14932 26630 14962 26682
rect 14962 26630 14974 26682
rect 14974 26630 14988 26682
rect 15012 26630 15026 26682
rect 15026 26630 15038 26682
rect 15038 26630 15068 26682
rect 15092 26630 15102 26682
rect 15102 26630 15148 26682
rect 14852 26628 14908 26630
rect 14932 26628 14988 26630
rect 15012 26628 15068 26630
rect 15092 26628 15148 26630
rect 14852 25594 14908 25596
rect 14932 25594 14988 25596
rect 15012 25594 15068 25596
rect 15092 25594 15148 25596
rect 14852 25542 14898 25594
rect 14898 25542 14908 25594
rect 14932 25542 14962 25594
rect 14962 25542 14974 25594
rect 14974 25542 14988 25594
rect 15012 25542 15026 25594
rect 15026 25542 15038 25594
rect 15038 25542 15068 25594
rect 15092 25542 15102 25594
rect 15102 25542 15148 25594
rect 14852 25540 14908 25542
rect 14932 25540 14988 25542
rect 15012 25540 15068 25542
rect 15092 25540 15148 25542
rect 10220 16346 10276 16348
rect 10300 16346 10356 16348
rect 10380 16346 10436 16348
rect 10460 16346 10516 16348
rect 10220 16294 10266 16346
rect 10266 16294 10276 16346
rect 10300 16294 10330 16346
rect 10330 16294 10342 16346
rect 10342 16294 10356 16346
rect 10380 16294 10394 16346
rect 10394 16294 10406 16346
rect 10406 16294 10436 16346
rect 10460 16294 10470 16346
rect 10470 16294 10516 16346
rect 10220 16292 10276 16294
rect 10300 16292 10356 16294
rect 10380 16292 10436 16294
rect 10460 16292 10516 16294
rect 10220 15258 10276 15260
rect 10300 15258 10356 15260
rect 10380 15258 10436 15260
rect 10460 15258 10516 15260
rect 10220 15206 10266 15258
rect 10266 15206 10276 15258
rect 10300 15206 10330 15258
rect 10330 15206 10342 15258
rect 10342 15206 10356 15258
rect 10380 15206 10394 15258
rect 10394 15206 10406 15258
rect 10406 15206 10436 15258
rect 10460 15206 10470 15258
rect 10470 15206 10516 15258
rect 10220 15204 10276 15206
rect 10300 15204 10356 15206
rect 10380 15204 10436 15206
rect 10460 15204 10516 15206
rect 10966 15408 11022 15464
rect 14852 24506 14908 24508
rect 14932 24506 14988 24508
rect 15012 24506 15068 24508
rect 15092 24506 15148 24508
rect 14852 24454 14898 24506
rect 14898 24454 14908 24506
rect 14932 24454 14962 24506
rect 14962 24454 14974 24506
rect 14974 24454 14988 24506
rect 15012 24454 15026 24506
rect 15026 24454 15038 24506
rect 15038 24454 15068 24506
rect 15092 24454 15102 24506
rect 15102 24454 15148 24506
rect 14852 24452 14908 24454
rect 14932 24452 14988 24454
rect 15012 24452 15068 24454
rect 15092 24452 15148 24454
rect 14852 23418 14908 23420
rect 14932 23418 14988 23420
rect 15012 23418 15068 23420
rect 15092 23418 15148 23420
rect 14852 23366 14898 23418
rect 14898 23366 14908 23418
rect 14932 23366 14962 23418
rect 14962 23366 14974 23418
rect 14974 23366 14988 23418
rect 15012 23366 15026 23418
rect 15026 23366 15038 23418
rect 15038 23366 15068 23418
rect 15092 23366 15102 23418
rect 15102 23366 15148 23418
rect 14852 23364 14908 23366
rect 14932 23364 14988 23366
rect 15012 23364 15068 23366
rect 15092 23364 15148 23366
rect 12714 17040 12770 17096
rect 10220 14170 10276 14172
rect 10300 14170 10356 14172
rect 10380 14170 10436 14172
rect 10460 14170 10516 14172
rect 10220 14118 10266 14170
rect 10266 14118 10276 14170
rect 10300 14118 10330 14170
rect 10330 14118 10342 14170
rect 10342 14118 10356 14170
rect 10380 14118 10394 14170
rect 10394 14118 10406 14170
rect 10406 14118 10436 14170
rect 10460 14118 10470 14170
rect 10470 14118 10516 14170
rect 10220 14116 10276 14118
rect 10300 14116 10356 14118
rect 10380 14116 10436 14118
rect 10460 14116 10516 14118
rect 9494 13676 9496 13696
rect 9496 13676 9548 13696
rect 9548 13676 9550 13696
rect 9494 13640 9550 13676
rect 7470 9560 7526 9616
rect 5588 9274 5644 9276
rect 5668 9274 5724 9276
rect 5748 9274 5804 9276
rect 5828 9274 5884 9276
rect 5588 9222 5634 9274
rect 5634 9222 5644 9274
rect 5668 9222 5698 9274
rect 5698 9222 5710 9274
rect 5710 9222 5724 9274
rect 5748 9222 5762 9274
rect 5762 9222 5774 9274
rect 5774 9222 5804 9274
rect 5828 9222 5838 9274
rect 5838 9222 5884 9274
rect 5588 9220 5644 9222
rect 5668 9220 5724 9222
rect 5748 9220 5804 9222
rect 5828 9220 5884 9222
rect 1858 8916 1860 8936
rect 1860 8916 1912 8936
rect 1912 8916 1914 8936
rect 1858 8880 1914 8916
rect 1766 8336 1822 8392
rect 1398 8200 1454 8256
rect 5588 8186 5644 8188
rect 5668 8186 5724 8188
rect 5748 8186 5804 8188
rect 5828 8186 5884 8188
rect 5588 8134 5634 8186
rect 5634 8134 5644 8186
rect 5668 8134 5698 8186
rect 5698 8134 5710 8186
rect 5710 8134 5724 8186
rect 5748 8134 5762 8186
rect 5762 8134 5774 8186
rect 5774 8134 5804 8186
rect 5828 8134 5838 8186
rect 5838 8134 5884 8186
rect 5588 8132 5644 8134
rect 5668 8132 5724 8134
rect 5748 8132 5804 8134
rect 5828 8132 5884 8134
rect 5588 7098 5644 7100
rect 5668 7098 5724 7100
rect 5748 7098 5804 7100
rect 5828 7098 5884 7100
rect 5588 7046 5634 7098
rect 5634 7046 5644 7098
rect 5668 7046 5698 7098
rect 5698 7046 5710 7098
rect 5710 7046 5724 7098
rect 5748 7046 5762 7098
rect 5762 7046 5774 7098
rect 5774 7046 5804 7098
rect 5828 7046 5838 7098
rect 5838 7046 5884 7098
rect 5588 7044 5644 7046
rect 5668 7044 5724 7046
rect 5748 7044 5804 7046
rect 5828 7044 5884 7046
rect 9126 9580 9182 9616
rect 9126 9560 9128 9580
rect 9128 9560 9180 9580
rect 9180 9560 9182 9580
rect 10220 13082 10276 13084
rect 10300 13082 10356 13084
rect 10380 13082 10436 13084
rect 10460 13082 10516 13084
rect 10220 13030 10266 13082
rect 10266 13030 10276 13082
rect 10300 13030 10330 13082
rect 10330 13030 10342 13082
rect 10342 13030 10356 13082
rect 10380 13030 10394 13082
rect 10394 13030 10406 13082
rect 10406 13030 10436 13082
rect 10460 13030 10470 13082
rect 10470 13030 10516 13082
rect 10220 13028 10276 13030
rect 10300 13028 10356 13030
rect 10380 13028 10436 13030
rect 10460 13028 10516 13030
rect 10220 11994 10276 11996
rect 10300 11994 10356 11996
rect 10380 11994 10436 11996
rect 10460 11994 10516 11996
rect 10220 11942 10266 11994
rect 10266 11942 10276 11994
rect 10300 11942 10330 11994
rect 10330 11942 10342 11994
rect 10342 11942 10356 11994
rect 10380 11942 10394 11994
rect 10394 11942 10406 11994
rect 10406 11942 10436 11994
rect 10460 11942 10470 11994
rect 10470 11942 10516 11994
rect 10220 11940 10276 11942
rect 10300 11940 10356 11942
rect 10380 11940 10436 11942
rect 10460 11940 10516 11942
rect 10230 11756 10286 11792
rect 10230 11736 10232 11756
rect 10232 11736 10284 11756
rect 10284 11736 10286 11756
rect 10322 11192 10378 11248
rect 10966 11736 11022 11792
rect 10220 10906 10276 10908
rect 10300 10906 10356 10908
rect 10380 10906 10436 10908
rect 10460 10906 10516 10908
rect 10220 10854 10266 10906
rect 10266 10854 10276 10906
rect 10300 10854 10330 10906
rect 10330 10854 10342 10906
rect 10342 10854 10356 10906
rect 10380 10854 10394 10906
rect 10394 10854 10406 10906
rect 10406 10854 10436 10906
rect 10460 10854 10470 10906
rect 10470 10854 10516 10906
rect 10220 10852 10276 10854
rect 10300 10852 10356 10854
rect 10380 10852 10436 10854
rect 10460 10852 10516 10854
rect 11150 11076 11206 11112
rect 11150 11056 11152 11076
rect 11152 11056 11204 11076
rect 11204 11056 11206 11076
rect 10220 9818 10276 9820
rect 10300 9818 10356 9820
rect 10380 9818 10436 9820
rect 10460 9818 10516 9820
rect 10220 9766 10266 9818
rect 10266 9766 10276 9818
rect 10300 9766 10330 9818
rect 10330 9766 10342 9818
rect 10342 9766 10356 9818
rect 10380 9766 10394 9818
rect 10394 9766 10406 9818
rect 10406 9766 10436 9818
rect 10460 9766 10470 9818
rect 10470 9766 10516 9818
rect 10220 9764 10276 9766
rect 10300 9764 10356 9766
rect 10380 9764 10436 9766
rect 10460 9764 10516 9766
rect 9678 8492 9734 8528
rect 9678 8472 9680 8492
rect 9680 8472 9732 8492
rect 9732 8472 9734 8492
rect 10220 8730 10276 8732
rect 10300 8730 10356 8732
rect 10380 8730 10436 8732
rect 10460 8730 10516 8732
rect 10220 8678 10266 8730
rect 10266 8678 10276 8730
rect 10300 8678 10330 8730
rect 10330 8678 10342 8730
rect 10342 8678 10356 8730
rect 10380 8678 10394 8730
rect 10394 8678 10406 8730
rect 10406 8678 10436 8730
rect 10460 8678 10470 8730
rect 10470 8678 10516 8730
rect 10220 8676 10276 8678
rect 10300 8676 10356 8678
rect 10380 8676 10436 8678
rect 10460 8676 10516 8678
rect 10046 7928 10102 7984
rect 5588 6010 5644 6012
rect 5668 6010 5724 6012
rect 5748 6010 5804 6012
rect 5828 6010 5884 6012
rect 5588 5958 5634 6010
rect 5634 5958 5644 6010
rect 5668 5958 5698 6010
rect 5698 5958 5710 6010
rect 5710 5958 5724 6010
rect 5748 5958 5762 6010
rect 5762 5958 5774 6010
rect 5774 5958 5804 6010
rect 5828 5958 5838 6010
rect 5838 5958 5884 6010
rect 5588 5956 5644 5958
rect 5668 5956 5724 5958
rect 5748 5956 5804 5958
rect 5828 5956 5884 5958
rect 8482 5908 8538 5944
rect 8482 5888 8484 5908
rect 8484 5888 8536 5908
rect 8536 5888 8538 5908
rect 1490 5516 1492 5536
rect 1492 5516 1544 5536
rect 1544 5516 1546 5536
rect 1490 5480 1546 5516
rect 5588 4922 5644 4924
rect 5668 4922 5724 4924
rect 5748 4922 5804 4924
rect 5828 4922 5884 4924
rect 5588 4870 5634 4922
rect 5634 4870 5644 4922
rect 5668 4870 5698 4922
rect 5698 4870 5710 4922
rect 5710 4870 5724 4922
rect 5748 4870 5762 4922
rect 5762 4870 5774 4922
rect 5774 4870 5804 4922
rect 5828 4870 5838 4922
rect 5838 4870 5884 4922
rect 5588 4868 5644 4870
rect 5668 4868 5724 4870
rect 5748 4868 5804 4870
rect 5828 4868 5884 4870
rect 10220 7642 10276 7644
rect 10300 7642 10356 7644
rect 10380 7642 10436 7644
rect 10460 7642 10516 7644
rect 10220 7590 10266 7642
rect 10266 7590 10276 7642
rect 10300 7590 10330 7642
rect 10330 7590 10342 7642
rect 10342 7590 10356 7642
rect 10380 7590 10394 7642
rect 10394 7590 10406 7642
rect 10406 7590 10436 7642
rect 10460 7590 10470 7642
rect 10470 7590 10516 7642
rect 10220 7588 10276 7590
rect 10300 7588 10356 7590
rect 10380 7588 10436 7590
rect 10460 7588 10516 7590
rect 10220 6554 10276 6556
rect 10300 6554 10356 6556
rect 10380 6554 10436 6556
rect 10460 6554 10516 6556
rect 10220 6502 10266 6554
rect 10266 6502 10276 6554
rect 10300 6502 10330 6554
rect 10330 6502 10342 6554
rect 10342 6502 10356 6554
rect 10380 6502 10394 6554
rect 10394 6502 10406 6554
rect 10406 6502 10436 6554
rect 10460 6502 10470 6554
rect 10470 6502 10516 6554
rect 10220 6500 10276 6502
rect 10300 6500 10356 6502
rect 10380 6500 10436 6502
rect 10460 6500 10516 6502
rect 10598 5652 10600 5672
rect 10600 5652 10652 5672
rect 10652 5652 10654 5672
rect 10598 5616 10654 5652
rect 10220 5466 10276 5468
rect 10300 5466 10356 5468
rect 10380 5466 10436 5468
rect 10460 5466 10516 5468
rect 10220 5414 10266 5466
rect 10266 5414 10276 5466
rect 10300 5414 10330 5466
rect 10330 5414 10342 5466
rect 10342 5414 10356 5466
rect 10380 5414 10394 5466
rect 10394 5414 10406 5466
rect 10406 5414 10436 5466
rect 10460 5414 10470 5466
rect 10470 5414 10516 5466
rect 10220 5412 10276 5414
rect 10300 5412 10356 5414
rect 10380 5412 10436 5414
rect 10460 5412 10516 5414
rect 5588 3834 5644 3836
rect 5668 3834 5724 3836
rect 5748 3834 5804 3836
rect 5828 3834 5884 3836
rect 5588 3782 5634 3834
rect 5634 3782 5644 3834
rect 5668 3782 5698 3834
rect 5698 3782 5710 3834
rect 5710 3782 5724 3834
rect 5748 3782 5762 3834
rect 5762 3782 5774 3834
rect 5774 3782 5804 3834
rect 5828 3782 5838 3834
rect 5838 3782 5884 3834
rect 5588 3780 5644 3782
rect 5668 3780 5724 3782
rect 5748 3780 5804 3782
rect 5828 3780 5884 3782
rect 10220 4378 10276 4380
rect 10300 4378 10356 4380
rect 10380 4378 10436 4380
rect 10460 4378 10516 4380
rect 10220 4326 10266 4378
rect 10266 4326 10276 4378
rect 10300 4326 10330 4378
rect 10330 4326 10342 4378
rect 10342 4326 10356 4378
rect 10380 4326 10394 4378
rect 10394 4326 10406 4378
rect 10406 4326 10436 4378
rect 10460 4326 10470 4378
rect 10470 4326 10516 4378
rect 10220 4324 10276 4326
rect 10300 4324 10356 4326
rect 10380 4324 10436 4326
rect 10460 4324 10516 4326
rect 12898 16396 12900 16416
rect 12900 16396 12952 16416
rect 12952 16396 12954 16416
rect 12898 16360 12954 16396
rect 13358 16532 13360 16552
rect 13360 16532 13412 16552
rect 13412 16532 13414 16552
rect 13358 16496 13414 16532
rect 14852 22330 14908 22332
rect 14932 22330 14988 22332
rect 15012 22330 15068 22332
rect 15092 22330 15148 22332
rect 14852 22278 14898 22330
rect 14898 22278 14908 22330
rect 14932 22278 14962 22330
rect 14962 22278 14974 22330
rect 14974 22278 14988 22330
rect 15012 22278 15026 22330
rect 15026 22278 15038 22330
rect 15038 22278 15068 22330
rect 15092 22278 15102 22330
rect 15102 22278 15148 22330
rect 14852 22276 14908 22278
rect 14932 22276 14988 22278
rect 15012 22276 15068 22278
rect 15092 22276 15148 22278
rect 14852 21242 14908 21244
rect 14932 21242 14988 21244
rect 15012 21242 15068 21244
rect 15092 21242 15148 21244
rect 14852 21190 14898 21242
rect 14898 21190 14908 21242
rect 14932 21190 14962 21242
rect 14962 21190 14974 21242
rect 14974 21190 14988 21242
rect 15012 21190 15026 21242
rect 15026 21190 15038 21242
rect 15038 21190 15068 21242
rect 15092 21190 15102 21242
rect 15102 21190 15148 21242
rect 14852 21188 14908 21190
rect 14932 21188 14988 21190
rect 15012 21188 15068 21190
rect 15092 21188 15148 21190
rect 13818 16632 13874 16688
rect 13542 16224 13598 16280
rect 14094 16632 14150 16688
rect 14002 16360 14058 16416
rect 14186 16360 14242 16416
rect 12990 15408 13046 15464
rect 14002 15544 14058 15600
rect 13266 14456 13322 14512
rect 13174 14320 13230 14376
rect 13174 13640 13230 13696
rect 14852 20154 14908 20156
rect 14932 20154 14988 20156
rect 15012 20154 15068 20156
rect 15092 20154 15148 20156
rect 14852 20102 14898 20154
rect 14898 20102 14908 20154
rect 14932 20102 14962 20154
rect 14962 20102 14974 20154
rect 14974 20102 14988 20154
rect 15012 20102 15026 20154
rect 15026 20102 15038 20154
rect 15038 20102 15068 20154
rect 15092 20102 15102 20154
rect 15102 20102 15148 20154
rect 14852 20100 14908 20102
rect 14932 20100 14988 20102
rect 15012 20100 15068 20102
rect 15092 20100 15148 20102
rect 14852 19066 14908 19068
rect 14932 19066 14988 19068
rect 15012 19066 15068 19068
rect 15092 19066 15148 19068
rect 14852 19014 14898 19066
rect 14898 19014 14908 19066
rect 14932 19014 14962 19066
rect 14962 19014 14974 19066
rect 14974 19014 14988 19066
rect 15012 19014 15026 19066
rect 15026 19014 15038 19066
rect 15038 19014 15068 19066
rect 15092 19014 15102 19066
rect 15102 19014 15148 19066
rect 14852 19012 14908 19014
rect 14932 19012 14988 19014
rect 15012 19012 15068 19014
rect 15092 19012 15148 19014
rect 14462 17040 14518 17096
rect 14370 16904 14426 16960
rect 14462 16632 14518 16688
rect 14278 14864 14334 14920
rect 14554 16108 14610 16144
rect 14554 16088 14556 16108
rect 14556 16088 14608 16108
rect 14608 16088 14610 16108
rect 14462 14884 14518 14920
rect 14462 14864 14464 14884
rect 14464 14864 14516 14884
rect 14516 14864 14518 14884
rect 13818 12180 13820 12200
rect 13820 12180 13872 12200
rect 13872 12180 13874 12200
rect 13818 12144 13874 12180
rect 12346 8472 12402 8528
rect 14852 17978 14908 17980
rect 14932 17978 14988 17980
rect 15012 17978 15068 17980
rect 15092 17978 15148 17980
rect 14852 17926 14898 17978
rect 14898 17926 14908 17978
rect 14932 17926 14962 17978
rect 14962 17926 14974 17978
rect 14974 17926 14988 17978
rect 15012 17926 15026 17978
rect 15026 17926 15038 17978
rect 15038 17926 15068 17978
rect 15092 17926 15102 17978
rect 15102 17926 15148 17978
rect 14852 17924 14908 17926
rect 14932 17924 14988 17926
rect 15012 17924 15068 17926
rect 15092 17924 15148 17926
rect 14852 16890 14908 16892
rect 14932 16890 14988 16892
rect 15012 16890 15068 16892
rect 15092 16890 15148 16892
rect 14852 16838 14898 16890
rect 14898 16838 14908 16890
rect 14932 16838 14962 16890
rect 14962 16838 14974 16890
rect 14974 16838 14988 16890
rect 15012 16838 15026 16890
rect 15026 16838 15038 16890
rect 15038 16838 15068 16890
rect 15092 16838 15102 16890
rect 15102 16838 15148 16890
rect 14852 16836 14908 16838
rect 14932 16836 14988 16838
rect 15012 16836 15068 16838
rect 15092 16836 15148 16838
rect 15198 16396 15200 16416
rect 15200 16396 15252 16416
rect 15252 16396 15254 16416
rect 15198 16360 15254 16396
rect 14852 15802 14908 15804
rect 14932 15802 14988 15804
rect 15012 15802 15068 15804
rect 15092 15802 15148 15804
rect 14852 15750 14898 15802
rect 14898 15750 14908 15802
rect 14932 15750 14962 15802
rect 14962 15750 14974 15802
rect 14974 15750 14988 15802
rect 15012 15750 15026 15802
rect 15026 15750 15038 15802
rect 15038 15750 15068 15802
rect 15092 15750 15102 15802
rect 15102 15750 15148 15802
rect 14852 15748 14908 15750
rect 14932 15748 14988 15750
rect 15012 15748 15068 15750
rect 15092 15748 15148 15750
rect 14852 14714 14908 14716
rect 14932 14714 14988 14716
rect 15012 14714 15068 14716
rect 15092 14714 15148 14716
rect 14852 14662 14898 14714
rect 14898 14662 14908 14714
rect 14932 14662 14962 14714
rect 14962 14662 14974 14714
rect 14974 14662 14988 14714
rect 15012 14662 15026 14714
rect 15026 14662 15038 14714
rect 15038 14662 15068 14714
rect 15092 14662 15102 14714
rect 15102 14662 15148 14714
rect 14852 14660 14908 14662
rect 14932 14660 14988 14662
rect 15012 14660 15068 14662
rect 15092 14660 15148 14662
rect 15198 14456 15254 14512
rect 14852 13626 14908 13628
rect 14932 13626 14988 13628
rect 15012 13626 15068 13628
rect 15092 13626 15148 13628
rect 14852 13574 14898 13626
rect 14898 13574 14908 13626
rect 14932 13574 14962 13626
rect 14962 13574 14974 13626
rect 14974 13574 14988 13626
rect 15012 13574 15026 13626
rect 15026 13574 15038 13626
rect 15038 13574 15068 13626
rect 15092 13574 15102 13626
rect 15102 13574 15148 13626
rect 14852 13572 14908 13574
rect 14932 13572 14988 13574
rect 15012 13572 15068 13574
rect 15092 13572 15148 13574
rect 14852 12538 14908 12540
rect 14932 12538 14988 12540
rect 15012 12538 15068 12540
rect 15092 12538 15148 12540
rect 14852 12486 14898 12538
rect 14898 12486 14908 12538
rect 14932 12486 14962 12538
rect 14962 12486 14974 12538
rect 14974 12486 14988 12538
rect 15012 12486 15026 12538
rect 15026 12486 15038 12538
rect 15038 12486 15068 12538
rect 15092 12486 15102 12538
rect 15102 12486 15148 12538
rect 14852 12484 14908 12486
rect 14932 12484 14988 12486
rect 15012 12484 15068 12486
rect 15092 12484 15148 12486
rect 14738 12280 14794 12336
rect 15382 16496 15438 16552
rect 15382 15972 15438 16008
rect 15382 15952 15384 15972
rect 15384 15952 15436 15972
rect 15436 15952 15438 15972
rect 15382 15544 15438 15600
rect 15198 11872 15254 11928
rect 14852 11450 14908 11452
rect 14932 11450 14988 11452
rect 15012 11450 15068 11452
rect 15092 11450 15148 11452
rect 14852 11398 14898 11450
rect 14898 11398 14908 11450
rect 14932 11398 14962 11450
rect 14962 11398 14974 11450
rect 14974 11398 14988 11450
rect 15012 11398 15026 11450
rect 15026 11398 15038 11450
rect 15038 11398 15068 11450
rect 15092 11398 15102 11450
rect 15102 11398 15148 11450
rect 14852 11396 14908 11398
rect 14932 11396 14988 11398
rect 15012 11396 15068 11398
rect 15092 11396 15148 11398
rect 8206 3440 8262 3496
rect 10220 3290 10276 3292
rect 10300 3290 10356 3292
rect 10380 3290 10436 3292
rect 10460 3290 10516 3292
rect 10220 3238 10266 3290
rect 10266 3238 10276 3290
rect 10300 3238 10330 3290
rect 10330 3238 10342 3290
rect 10342 3238 10356 3290
rect 10380 3238 10394 3290
rect 10394 3238 10406 3290
rect 10406 3238 10436 3290
rect 10460 3238 10470 3290
rect 10470 3238 10516 3290
rect 10220 3236 10276 3238
rect 10300 3236 10356 3238
rect 10380 3236 10436 3238
rect 10460 3236 10516 3238
rect 12254 5072 12310 5128
rect 12530 4936 12586 4992
rect 15014 11212 15070 11248
rect 15014 11192 15016 11212
rect 15016 11192 15068 11212
rect 15068 11192 15070 11212
rect 17222 21292 17224 21312
rect 17224 21292 17276 21312
rect 17276 21292 17278 21312
rect 17222 21256 17278 21292
rect 19484 27226 19540 27228
rect 19564 27226 19620 27228
rect 19644 27226 19700 27228
rect 19724 27226 19780 27228
rect 19484 27174 19530 27226
rect 19530 27174 19540 27226
rect 19564 27174 19594 27226
rect 19594 27174 19606 27226
rect 19606 27174 19620 27226
rect 19644 27174 19658 27226
rect 19658 27174 19670 27226
rect 19670 27174 19700 27226
rect 19724 27174 19734 27226
rect 19734 27174 19780 27226
rect 19484 27172 19540 27174
rect 19564 27172 19620 27174
rect 19644 27172 19700 27174
rect 19724 27172 19780 27174
rect 19484 26138 19540 26140
rect 19564 26138 19620 26140
rect 19644 26138 19700 26140
rect 19724 26138 19780 26140
rect 19484 26086 19530 26138
rect 19530 26086 19540 26138
rect 19564 26086 19594 26138
rect 19594 26086 19606 26138
rect 19606 26086 19620 26138
rect 19644 26086 19658 26138
rect 19658 26086 19670 26138
rect 19670 26086 19700 26138
rect 19724 26086 19734 26138
rect 19734 26086 19780 26138
rect 19484 26084 19540 26086
rect 19564 26084 19620 26086
rect 19644 26084 19700 26086
rect 19724 26084 19780 26086
rect 19484 25050 19540 25052
rect 19564 25050 19620 25052
rect 19644 25050 19700 25052
rect 19724 25050 19780 25052
rect 19484 24998 19530 25050
rect 19530 24998 19540 25050
rect 19564 24998 19594 25050
rect 19594 24998 19606 25050
rect 19606 24998 19620 25050
rect 19644 24998 19658 25050
rect 19658 24998 19670 25050
rect 19670 24998 19700 25050
rect 19724 24998 19734 25050
rect 19734 24998 19780 25050
rect 19484 24996 19540 24998
rect 19564 24996 19620 24998
rect 19644 24996 19700 24998
rect 19724 24996 19780 24998
rect 19484 23962 19540 23964
rect 19564 23962 19620 23964
rect 19644 23962 19700 23964
rect 19724 23962 19780 23964
rect 19484 23910 19530 23962
rect 19530 23910 19540 23962
rect 19564 23910 19594 23962
rect 19594 23910 19606 23962
rect 19606 23910 19620 23962
rect 19644 23910 19658 23962
rect 19658 23910 19670 23962
rect 19670 23910 19700 23962
rect 19724 23910 19734 23962
rect 19734 23910 19780 23962
rect 19484 23908 19540 23910
rect 19564 23908 19620 23910
rect 19644 23908 19700 23910
rect 19724 23908 19780 23910
rect 19484 22874 19540 22876
rect 19564 22874 19620 22876
rect 19644 22874 19700 22876
rect 19724 22874 19780 22876
rect 19484 22822 19530 22874
rect 19530 22822 19540 22874
rect 19564 22822 19594 22874
rect 19594 22822 19606 22874
rect 19606 22822 19620 22874
rect 19644 22822 19658 22874
rect 19658 22822 19670 22874
rect 19670 22822 19700 22874
rect 19724 22822 19734 22874
rect 19734 22822 19780 22874
rect 19484 22820 19540 22822
rect 19564 22820 19620 22822
rect 19644 22820 19700 22822
rect 19724 22820 19780 22822
rect 19484 21786 19540 21788
rect 19564 21786 19620 21788
rect 19644 21786 19700 21788
rect 19724 21786 19780 21788
rect 19484 21734 19530 21786
rect 19530 21734 19540 21786
rect 19564 21734 19594 21786
rect 19594 21734 19606 21786
rect 19606 21734 19620 21786
rect 19644 21734 19658 21786
rect 19658 21734 19670 21786
rect 19670 21734 19700 21786
rect 19724 21734 19734 21786
rect 19734 21734 19780 21786
rect 19484 21732 19540 21734
rect 19564 21732 19620 21734
rect 19644 21732 19700 21734
rect 19724 21732 19780 21734
rect 19338 21256 19394 21312
rect 16486 17604 16542 17640
rect 16486 17584 16488 17604
rect 16488 17584 16540 17604
rect 16540 17584 16542 17604
rect 16210 15020 16266 15056
rect 16210 15000 16212 15020
rect 16212 15000 16264 15020
rect 16264 15000 16266 15020
rect 17130 15408 17186 15464
rect 16946 15000 17002 15056
rect 14852 10362 14908 10364
rect 14932 10362 14988 10364
rect 15012 10362 15068 10364
rect 15092 10362 15148 10364
rect 14852 10310 14898 10362
rect 14898 10310 14908 10362
rect 14932 10310 14962 10362
rect 14962 10310 14974 10362
rect 14974 10310 14988 10362
rect 15012 10310 15026 10362
rect 15026 10310 15038 10362
rect 15038 10310 15068 10362
rect 15092 10310 15102 10362
rect 15102 10310 15148 10362
rect 14852 10308 14908 10310
rect 14932 10308 14988 10310
rect 15012 10308 15068 10310
rect 15092 10308 15148 10310
rect 14852 9274 14908 9276
rect 14932 9274 14988 9276
rect 15012 9274 15068 9276
rect 15092 9274 15148 9276
rect 14852 9222 14898 9274
rect 14898 9222 14908 9274
rect 14932 9222 14962 9274
rect 14962 9222 14974 9274
rect 14974 9222 14988 9274
rect 15012 9222 15026 9274
rect 15026 9222 15038 9274
rect 15038 9222 15068 9274
rect 15092 9222 15102 9274
rect 15102 9222 15148 9274
rect 14852 9220 14908 9222
rect 14932 9220 14988 9222
rect 15012 9220 15068 9222
rect 15092 9220 15148 9222
rect 14852 8186 14908 8188
rect 14932 8186 14988 8188
rect 15012 8186 15068 8188
rect 15092 8186 15148 8188
rect 14852 8134 14898 8186
rect 14898 8134 14908 8186
rect 14932 8134 14962 8186
rect 14962 8134 14974 8186
rect 14974 8134 14988 8186
rect 15012 8134 15026 8186
rect 15026 8134 15038 8186
rect 15038 8134 15068 8186
rect 15092 8134 15102 8186
rect 15102 8134 15148 8186
rect 14852 8132 14908 8134
rect 14932 8132 14988 8134
rect 15012 8132 15068 8134
rect 15092 8132 15148 8134
rect 14852 7098 14908 7100
rect 14932 7098 14988 7100
rect 15012 7098 15068 7100
rect 15092 7098 15148 7100
rect 14852 7046 14898 7098
rect 14898 7046 14908 7098
rect 14932 7046 14962 7098
rect 14962 7046 14974 7098
rect 14974 7046 14988 7098
rect 15012 7046 15026 7098
rect 15026 7046 15038 7098
rect 15038 7046 15068 7098
rect 15092 7046 15102 7098
rect 15102 7046 15148 7098
rect 14852 7044 14908 7046
rect 14932 7044 14988 7046
rect 15012 7044 15068 7046
rect 15092 7044 15148 7046
rect 14852 6010 14908 6012
rect 14932 6010 14988 6012
rect 15012 6010 15068 6012
rect 15092 6010 15148 6012
rect 14852 5958 14898 6010
rect 14898 5958 14908 6010
rect 14932 5958 14962 6010
rect 14962 5958 14974 6010
rect 14974 5958 14988 6010
rect 15012 5958 15026 6010
rect 15026 5958 15038 6010
rect 15038 5958 15068 6010
rect 15092 5958 15102 6010
rect 15102 5958 15148 6010
rect 14852 5956 14908 5958
rect 14932 5956 14988 5958
rect 15012 5956 15068 5958
rect 15092 5956 15148 5958
rect 14852 4922 14908 4924
rect 14932 4922 14988 4924
rect 15012 4922 15068 4924
rect 15092 4922 15148 4924
rect 14852 4870 14898 4922
rect 14898 4870 14908 4922
rect 14932 4870 14962 4922
rect 14962 4870 14974 4922
rect 14974 4870 14988 4922
rect 15012 4870 15026 4922
rect 15026 4870 15038 4922
rect 15038 4870 15068 4922
rect 15092 4870 15102 4922
rect 15102 4870 15148 4922
rect 14852 4868 14908 4870
rect 14932 4868 14988 4870
rect 15012 4868 15068 4870
rect 15092 4868 15148 4870
rect 14852 3834 14908 3836
rect 14932 3834 14988 3836
rect 15012 3834 15068 3836
rect 15092 3834 15148 3836
rect 14852 3782 14898 3834
rect 14898 3782 14908 3834
rect 14932 3782 14962 3834
rect 14962 3782 14974 3834
rect 14974 3782 14988 3834
rect 15012 3782 15026 3834
rect 15026 3782 15038 3834
rect 15038 3782 15068 3834
rect 15092 3782 15102 3834
rect 15102 3782 15148 3834
rect 14852 3780 14908 3782
rect 14932 3780 14988 3782
rect 15012 3780 15068 3782
rect 15092 3780 15148 3782
rect 5588 2746 5644 2748
rect 5668 2746 5724 2748
rect 5748 2746 5804 2748
rect 5828 2746 5884 2748
rect 5588 2694 5634 2746
rect 5634 2694 5644 2746
rect 5668 2694 5698 2746
rect 5698 2694 5710 2746
rect 5710 2694 5724 2746
rect 5748 2694 5762 2746
rect 5762 2694 5774 2746
rect 5774 2694 5804 2746
rect 5828 2694 5838 2746
rect 5838 2694 5884 2746
rect 5588 2692 5644 2694
rect 5668 2692 5724 2694
rect 5748 2692 5804 2694
rect 5828 2692 5884 2694
rect 14852 2746 14908 2748
rect 14932 2746 14988 2748
rect 15012 2746 15068 2748
rect 15092 2746 15148 2748
rect 14852 2694 14898 2746
rect 14898 2694 14908 2746
rect 14932 2694 14962 2746
rect 14962 2694 14974 2746
rect 14974 2694 14988 2746
rect 15012 2694 15026 2746
rect 15026 2694 15038 2746
rect 15038 2694 15068 2746
rect 15092 2694 15102 2746
rect 15102 2694 15148 2746
rect 14852 2692 14908 2694
rect 14932 2692 14988 2694
rect 15012 2692 15068 2694
rect 15092 2692 15148 2694
rect 2226 2080 2282 2136
rect 10220 2202 10276 2204
rect 10300 2202 10356 2204
rect 10380 2202 10436 2204
rect 10460 2202 10516 2204
rect 10220 2150 10266 2202
rect 10266 2150 10276 2202
rect 10300 2150 10330 2202
rect 10330 2150 10342 2202
rect 10342 2150 10356 2202
rect 10380 2150 10394 2202
rect 10394 2150 10406 2202
rect 10406 2150 10436 2202
rect 10460 2150 10470 2202
rect 10470 2150 10516 2202
rect 10220 2148 10276 2150
rect 10300 2148 10356 2150
rect 10380 2148 10436 2150
rect 10460 2148 10516 2150
rect 17038 14356 17040 14376
rect 17040 14356 17092 14376
rect 17092 14356 17094 14376
rect 17038 14320 17094 14356
rect 19484 20698 19540 20700
rect 19564 20698 19620 20700
rect 19644 20698 19700 20700
rect 19724 20698 19780 20700
rect 19484 20646 19530 20698
rect 19530 20646 19540 20698
rect 19564 20646 19594 20698
rect 19594 20646 19606 20698
rect 19606 20646 19620 20698
rect 19644 20646 19658 20698
rect 19658 20646 19670 20698
rect 19670 20646 19700 20698
rect 19724 20646 19734 20698
rect 19734 20646 19780 20698
rect 19484 20644 19540 20646
rect 19564 20644 19620 20646
rect 19644 20644 19700 20646
rect 19724 20644 19780 20646
rect 19484 19610 19540 19612
rect 19564 19610 19620 19612
rect 19644 19610 19700 19612
rect 19724 19610 19780 19612
rect 19484 19558 19530 19610
rect 19530 19558 19540 19610
rect 19564 19558 19594 19610
rect 19594 19558 19606 19610
rect 19606 19558 19620 19610
rect 19644 19558 19658 19610
rect 19658 19558 19670 19610
rect 19670 19558 19700 19610
rect 19724 19558 19734 19610
rect 19734 19558 19780 19610
rect 19484 19556 19540 19558
rect 19564 19556 19620 19558
rect 19644 19556 19700 19558
rect 19724 19556 19780 19558
rect 19484 18522 19540 18524
rect 19564 18522 19620 18524
rect 19644 18522 19700 18524
rect 19724 18522 19780 18524
rect 19484 18470 19530 18522
rect 19530 18470 19540 18522
rect 19564 18470 19594 18522
rect 19594 18470 19606 18522
rect 19606 18470 19620 18522
rect 19644 18470 19658 18522
rect 19658 18470 19670 18522
rect 19670 18470 19700 18522
rect 19724 18470 19734 18522
rect 19734 18470 19780 18522
rect 19484 18468 19540 18470
rect 19564 18468 19620 18470
rect 19644 18468 19700 18470
rect 19724 18468 19780 18470
rect 18326 17176 18382 17232
rect 17682 15000 17738 15056
rect 17866 15000 17922 15056
rect 17590 13368 17646 13424
rect 17498 12008 17554 12064
rect 16118 8880 16174 8936
rect 16578 5652 16580 5672
rect 16580 5652 16632 5672
rect 16632 5652 16634 5672
rect 16578 5616 16634 5652
rect 19484 17434 19540 17436
rect 19564 17434 19620 17436
rect 19644 17434 19700 17436
rect 19724 17434 19780 17436
rect 19484 17382 19530 17434
rect 19530 17382 19540 17434
rect 19564 17382 19594 17434
rect 19594 17382 19606 17434
rect 19606 17382 19620 17434
rect 19644 17382 19658 17434
rect 19658 17382 19670 17434
rect 19670 17382 19700 17434
rect 19724 17382 19734 17434
rect 19734 17382 19780 17434
rect 19484 17380 19540 17382
rect 19564 17380 19620 17382
rect 19644 17380 19700 17382
rect 19724 17380 19780 17382
rect 18234 12144 18290 12200
rect 19484 16346 19540 16348
rect 19564 16346 19620 16348
rect 19644 16346 19700 16348
rect 19724 16346 19780 16348
rect 19484 16294 19530 16346
rect 19530 16294 19540 16346
rect 19564 16294 19594 16346
rect 19594 16294 19606 16346
rect 19606 16294 19620 16346
rect 19644 16294 19658 16346
rect 19658 16294 19670 16346
rect 19670 16294 19700 16346
rect 19724 16294 19734 16346
rect 19734 16294 19780 16346
rect 19484 16292 19540 16294
rect 19564 16292 19620 16294
rect 19644 16292 19700 16294
rect 19724 16292 19780 16294
rect 19338 16244 19394 16280
rect 19338 16224 19340 16244
rect 19340 16224 19392 16244
rect 19392 16224 19394 16244
rect 19484 15258 19540 15260
rect 19564 15258 19620 15260
rect 19644 15258 19700 15260
rect 19724 15258 19780 15260
rect 19484 15206 19530 15258
rect 19530 15206 19540 15258
rect 19564 15206 19594 15258
rect 19594 15206 19606 15258
rect 19606 15206 19620 15258
rect 19644 15206 19658 15258
rect 19658 15206 19670 15258
rect 19670 15206 19700 15258
rect 19724 15206 19734 15258
rect 19734 15206 19780 15258
rect 19484 15204 19540 15206
rect 19564 15204 19620 15206
rect 19644 15204 19700 15206
rect 19724 15204 19780 15206
rect 19798 15036 19800 15056
rect 19800 15036 19852 15056
rect 19852 15036 19854 15056
rect 19798 15000 19854 15036
rect 21086 19660 21088 19680
rect 21088 19660 21140 19680
rect 21140 19660 21142 19680
rect 21086 19624 21142 19660
rect 24116 26682 24172 26684
rect 24196 26682 24252 26684
rect 24276 26682 24332 26684
rect 24356 26682 24412 26684
rect 24116 26630 24162 26682
rect 24162 26630 24172 26682
rect 24196 26630 24226 26682
rect 24226 26630 24238 26682
rect 24238 26630 24252 26682
rect 24276 26630 24290 26682
rect 24290 26630 24302 26682
rect 24302 26630 24332 26682
rect 24356 26630 24366 26682
rect 24366 26630 24412 26682
rect 24116 26628 24172 26630
rect 24196 26628 24252 26630
rect 24276 26628 24332 26630
rect 24356 26628 24412 26630
rect 19484 14170 19540 14172
rect 19564 14170 19620 14172
rect 19644 14170 19700 14172
rect 19724 14170 19780 14172
rect 19484 14118 19530 14170
rect 19530 14118 19540 14170
rect 19564 14118 19594 14170
rect 19594 14118 19606 14170
rect 19606 14118 19620 14170
rect 19644 14118 19658 14170
rect 19658 14118 19670 14170
rect 19670 14118 19700 14170
rect 19724 14118 19734 14170
rect 19734 14118 19780 14170
rect 19484 14116 19540 14118
rect 19564 14116 19620 14118
rect 19644 14116 19700 14118
rect 19724 14116 19780 14118
rect 19484 13082 19540 13084
rect 19564 13082 19620 13084
rect 19644 13082 19700 13084
rect 19724 13082 19780 13084
rect 19484 13030 19530 13082
rect 19530 13030 19540 13082
rect 19564 13030 19594 13082
rect 19594 13030 19606 13082
rect 19606 13030 19620 13082
rect 19644 13030 19658 13082
rect 19658 13030 19670 13082
rect 19670 13030 19700 13082
rect 19724 13030 19734 13082
rect 19734 13030 19780 13082
rect 19484 13028 19540 13030
rect 19564 13028 19620 13030
rect 19644 13028 19700 13030
rect 19724 13028 19780 13030
rect 19484 11994 19540 11996
rect 19564 11994 19620 11996
rect 19644 11994 19700 11996
rect 19724 11994 19780 11996
rect 19484 11942 19530 11994
rect 19530 11942 19540 11994
rect 19564 11942 19594 11994
rect 19594 11942 19606 11994
rect 19606 11942 19620 11994
rect 19644 11942 19658 11994
rect 19658 11942 19670 11994
rect 19670 11942 19700 11994
rect 19724 11942 19734 11994
rect 19734 11942 19780 11994
rect 19484 11940 19540 11942
rect 19564 11940 19620 11942
rect 19644 11940 19700 11942
rect 19724 11940 19780 11942
rect 19484 10906 19540 10908
rect 19564 10906 19620 10908
rect 19644 10906 19700 10908
rect 19724 10906 19780 10908
rect 19484 10854 19530 10906
rect 19530 10854 19540 10906
rect 19564 10854 19594 10906
rect 19594 10854 19606 10906
rect 19606 10854 19620 10906
rect 19644 10854 19658 10906
rect 19658 10854 19670 10906
rect 19670 10854 19700 10906
rect 19724 10854 19734 10906
rect 19734 10854 19780 10906
rect 19484 10852 19540 10854
rect 19564 10852 19620 10854
rect 19644 10852 19700 10854
rect 19724 10852 19780 10854
rect 19484 9818 19540 9820
rect 19564 9818 19620 9820
rect 19644 9818 19700 9820
rect 19724 9818 19780 9820
rect 19484 9766 19530 9818
rect 19530 9766 19540 9818
rect 19564 9766 19594 9818
rect 19594 9766 19606 9818
rect 19606 9766 19620 9818
rect 19644 9766 19658 9818
rect 19658 9766 19670 9818
rect 19670 9766 19700 9818
rect 19724 9766 19734 9818
rect 19734 9766 19780 9818
rect 19484 9764 19540 9766
rect 19564 9764 19620 9766
rect 19644 9764 19700 9766
rect 19724 9764 19780 9766
rect 19484 8730 19540 8732
rect 19564 8730 19620 8732
rect 19644 8730 19700 8732
rect 19724 8730 19780 8732
rect 19484 8678 19530 8730
rect 19530 8678 19540 8730
rect 19564 8678 19594 8730
rect 19594 8678 19606 8730
rect 19606 8678 19620 8730
rect 19644 8678 19658 8730
rect 19658 8678 19670 8730
rect 19670 8678 19700 8730
rect 19724 8678 19734 8730
rect 19734 8678 19780 8730
rect 19484 8676 19540 8678
rect 19564 8676 19620 8678
rect 19644 8676 19700 8678
rect 19724 8676 19780 8678
rect 18694 8356 18750 8392
rect 18694 8336 18696 8356
rect 18696 8336 18748 8356
rect 18748 8336 18750 8356
rect 19484 7642 19540 7644
rect 19564 7642 19620 7644
rect 19644 7642 19700 7644
rect 19724 7642 19780 7644
rect 19484 7590 19530 7642
rect 19530 7590 19540 7642
rect 19564 7590 19594 7642
rect 19594 7590 19606 7642
rect 19606 7590 19620 7642
rect 19644 7590 19658 7642
rect 19658 7590 19670 7642
rect 19670 7590 19700 7642
rect 19724 7590 19734 7642
rect 19734 7590 19780 7642
rect 19484 7588 19540 7590
rect 19564 7588 19620 7590
rect 19644 7588 19700 7590
rect 19724 7588 19780 7590
rect 19484 6554 19540 6556
rect 19564 6554 19620 6556
rect 19644 6554 19700 6556
rect 19724 6554 19780 6556
rect 19484 6502 19530 6554
rect 19530 6502 19540 6554
rect 19564 6502 19594 6554
rect 19594 6502 19606 6554
rect 19606 6502 19620 6554
rect 19644 6502 19658 6554
rect 19658 6502 19670 6554
rect 19670 6502 19700 6554
rect 19724 6502 19734 6554
rect 19734 6502 19780 6554
rect 19484 6500 19540 6502
rect 19564 6500 19620 6502
rect 19644 6500 19700 6502
rect 19724 6500 19780 6502
rect 19484 5466 19540 5468
rect 19564 5466 19620 5468
rect 19644 5466 19700 5468
rect 19724 5466 19780 5468
rect 19484 5414 19530 5466
rect 19530 5414 19540 5466
rect 19564 5414 19594 5466
rect 19594 5414 19606 5466
rect 19606 5414 19620 5466
rect 19644 5414 19658 5466
rect 19658 5414 19670 5466
rect 19670 5414 19700 5466
rect 19724 5414 19734 5466
rect 19734 5414 19780 5466
rect 19484 5412 19540 5414
rect 19564 5412 19620 5414
rect 19644 5412 19700 5414
rect 19724 5412 19780 5414
rect 19484 4378 19540 4380
rect 19564 4378 19620 4380
rect 19644 4378 19700 4380
rect 19724 4378 19780 4380
rect 19484 4326 19530 4378
rect 19530 4326 19540 4378
rect 19564 4326 19594 4378
rect 19594 4326 19606 4378
rect 19606 4326 19620 4378
rect 19644 4326 19658 4378
rect 19658 4326 19670 4378
rect 19670 4326 19700 4378
rect 19724 4326 19734 4378
rect 19734 4326 19780 4378
rect 19484 4324 19540 4326
rect 19564 4324 19620 4326
rect 19644 4324 19700 4326
rect 19724 4324 19780 4326
rect 19484 3290 19540 3292
rect 19564 3290 19620 3292
rect 19644 3290 19700 3292
rect 19724 3290 19780 3292
rect 19484 3238 19530 3290
rect 19530 3238 19540 3290
rect 19564 3238 19594 3290
rect 19594 3238 19606 3290
rect 19606 3238 19620 3290
rect 19644 3238 19658 3290
rect 19658 3238 19670 3290
rect 19670 3238 19700 3290
rect 19724 3238 19734 3290
rect 19734 3238 19780 3290
rect 19484 3236 19540 3238
rect 19564 3236 19620 3238
rect 19644 3236 19700 3238
rect 19724 3236 19780 3238
rect 20994 16088 21050 16144
rect 20442 15156 20498 15192
rect 20442 15136 20444 15156
rect 20444 15136 20496 15156
rect 20496 15136 20498 15156
rect 20718 15020 20774 15056
rect 20718 15000 20720 15020
rect 20720 15000 20772 15020
rect 20772 15000 20774 15020
rect 20810 12280 20866 12336
rect 22098 17584 22154 17640
rect 22098 15972 22154 16008
rect 22098 15952 22100 15972
rect 22100 15952 22152 15972
rect 22152 15952 22154 15972
rect 22006 15408 22062 15464
rect 22466 13268 22468 13288
rect 22468 13268 22520 13288
rect 22520 13268 22522 13288
rect 22466 13232 22522 13268
rect 22558 12164 22614 12200
rect 22558 12144 22560 12164
rect 22560 12144 22612 12164
rect 22612 12144 22614 12164
rect 24116 25594 24172 25596
rect 24196 25594 24252 25596
rect 24276 25594 24332 25596
rect 24356 25594 24412 25596
rect 24116 25542 24162 25594
rect 24162 25542 24172 25594
rect 24196 25542 24226 25594
rect 24226 25542 24238 25594
rect 24238 25542 24252 25594
rect 24276 25542 24290 25594
rect 24290 25542 24302 25594
rect 24302 25542 24332 25594
rect 24356 25542 24366 25594
rect 24366 25542 24412 25594
rect 24116 25540 24172 25542
rect 24196 25540 24252 25542
rect 24276 25540 24332 25542
rect 24356 25540 24412 25542
rect 24116 24506 24172 24508
rect 24196 24506 24252 24508
rect 24276 24506 24332 24508
rect 24356 24506 24412 24508
rect 24116 24454 24162 24506
rect 24162 24454 24172 24506
rect 24196 24454 24226 24506
rect 24226 24454 24238 24506
rect 24238 24454 24252 24506
rect 24276 24454 24290 24506
rect 24290 24454 24302 24506
rect 24302 24454 24332 24506
rect 24356 24454 24366 24506
rect 24366 24454 24412 24506
rect 24116 24452 24172 24454
rect 24196 24452 24252 24454
rect 24276 24452 24332 24454
rect 24356 24452 24412 24454
rect 24116 23418 24172 23420
rect 24196 23418 24252 23420
rect 24276 23418 24332 23420
rect 24356 23418 24412 23420
rect 24116 23366 24162 23418
rect 24162 23366 24172 23418
rect 24196 23366 24226 23418
rect 24226 23366 24238 23418
rect 24238 23366 24252 23418
rect 24276 23366 24290 23418
rect 24290 23366 24302 23418
rect 24302 23366 24332 23418
rect 24356 23366 24366 23418
rect 24366 23366 24412 23418
rect 24116 23364 24172 23366
rect 24196 23364 24252 23366
rect 24276 23364 24332 23366
rect 24356 23364 24412 23366
rect 24116 22330 24172 22332
rect 24196 22330 24252 22332
rect 24276 22330 24332 22332
rect 24356 22330 24412 22332
rect 24116 22278 24162 22330
rect 24162 22278 24172 22330
rect 24196 22278 24226 22330
rect 24226 22278 24238 22330
rect 24238 22278 24252 22330
rect 24276 22278 24290 22330
rect 24290 22278 24302 22330
rect 24302 22278 24332 22330
rect 24356 22278 24366 22330
rect 24366 22278 24412 22330
rect 24116 22276 24172 22278
rect 24196 22276 24252 22278
rect 24276 22276 24332 22278
rect 24356 22276 24412 22278
rect 28262 27920 28318 27976
rect 24116 21242 24172 21244
rect 24196 21242 24252 21244
rect 24276 21242 24332 21244
rect 24356 21242 24412 21244
rect 24116 21190 24162 21242
rect 24162 21190 24172 21242
rect 24196 21190 24226 21242
rect 24226 21190 24238 21242
rect 24238 21190 24252 21242
rect 24276 21190 24290 21242
rect 24290 21190 24302 21242
rect 24302 21190 24332 21242
rect 24356 21190 24366 21242
rect 24366 21190 24412 21242
rect 24116 21188 24172 21190
rect 24196 21188 24252 21190
rect 24276 21188 24332 21190
rect 24356 21188 24412 21190
rect 24116 20154 24172 20156
rect 24196 20154 24252 20156
rect 24276 20154 24332 20156
rect 24356 20154 24412 20156
rect 24116 20102 24162 20154
rect 24162 20102 24172 20154
rect 24196 20102 24226 20154
rect 24226 20102 24238 20154
rect 24238 20102 24252 20154
rect 24276 20102 24290 20154
rect 24290 20102 24302 20154
rect 24302 20102 24332 20154
rect 24356 20102 24366 20154
rect 24366 20102 24412 20154
rect 24116 20100 24172 20102
rect 24196 20100 24252 20102
rect 24276 20100 24332 20102
rect 24356 20100 24412 20102
rect 24116 19066 24172 19068
rect 24196 19066 24252 19068
rect 24276 19066 24332 19068
rect 24356 19066 24412 19068
rect 24116 19014 24162 19066
rect 24162 19014 24172 19066
rect 24196 19014 24226 19066
rect 24226 19014 24238 19066
rect 24238 19014 24252 19066
rect 24276 19014 24290 19066
rect 24290 19014 24302 19066
rect 24302 19014 24332 19066
rect 24356 19014 24366 19066
rect 24366 19014 24412 19066
rect 24116 19012 24172 19014
rect 24196 19012 24252 19014
rect 24276 19012 24332 19014
rect 24356 19012 24412 19014
rect 24116 17978 24172 17980
rect 24196 17978 24252 17980
rect 24276 17978 24332 17980
rect 24356 17978 24412 17980
rect 24116 17926 24162 17978
rect 24162 17926 24172 17978
rect 24196 17926 24226 17978
rect 24226 17926 24238 17978
rect 24238 17926 24252 17978
rect 24276 17926 24290 17978
rect 24290 17926 24302 17978
rect 24302 17926 24332 17978
rect 24356 17926 24366 17978
rect 24366 17926 24412 17978
rect 24116 17924 24172 17926
rect 24196 17924 24252 17926
rect 24276 17924 24332 17926
rect 24356 17924 24412 17926
rect 24116 16890 24172 16892
rect 24196 16890 24252 16892
rect 24276 16890 24332 16892
rect 24356 16890 24412 16892
rect 24116 16838 24162 16890
rect 24162 16838 24172 16890
rect 24196 16838 24226 16890
rect 24226 16838 24238 16890
rect 24238 16838 24252 16890
rect 24276 16838 24290 16890
rect 24290 16838 24302 16890
rect 24302 16838 24332 16890
rect 24356 16838 24366 16890
rect 24366 16838 24412 16890
rect 24116 16836 24172 16838
rect 24196 16836 24252 16838
rect 24276 16836 24332 16838
rect 24356 16836 24412 16838
rect 28354 26580 28410 26616
rect 28354 26560 28356 26580
rect 28356 26560 28408 26580
rect 28408 26560 28410 26580
rect 28354 25236 28356 25256
rect 28356 25236 28408 25256
rect 28408 25236 28410 25256
rect 28354 25200 28410 25236
rect 24116 15802 24172 15804
rect 24196 15802 24252 15804
rect 24276 15802 24332 15804
rect 24356 15802 24412 15804
rect 24116 15750 24162 15802
rect 24162 15750 24172 15802
rect 24196 15750 24226 15802
rect 24226 15750 24238 15802
rect 24238 15750 24252 15802
rect 24276 15750 24290 15802
rect 24290 15750 24302 15802
rect 24302 15750 24332 15802
rect 24356 15750 24366 15802
rect 24366 15750 24412 15802
rect 24116 15748 24172 15750
rect 24196 15748 24252 15750
rect 24276 15748 24332 15750
rect 24356 15748 24412 15750
rect 23846 15136 23902 15192
rect 23478 14864 23534 14920
rect 24116 14714 24172 14716
rect 24196 14714 24252 14716
rect 24276 14714 24332 14716
rect 24356 14714 24412 14716
rect 24116 14662 24162 14714
rect 24162 14662 24172 14714
rect 24196 14662 24226 14714
rect 24226 14662 24238 14714
rect 24238 14662 24252 14714
rect 24276 14662 24290 14714
rect 24290 14662 24302 14714
rect 24302 14662 24332 14714
rect 24356 14662 24366 14714
rect 24366 14662 24412 14714
rect 24116 14660 24172 14662
rect 24196 14660 24252 14662
rect 24276 14660 24332 14662
rect 24356 14660 24412 14662
rect 24116 13626 24172 13628
rect 24196 13626 24252 13628
rect 24276 13626 24332 13628
rect 24356 13626 24412 13628
rect 24116 13574 24162 13626
rect 24162 13574 24172 13626
rect 24196 13574 24226 13626
rect 24226 13574 24238 13626
rect 24238 13574 24252 13626
rect 24276 13574 24290 13626
rect 24290 13574 24302 13626
rect 24302 13574 24332 13626
rect 24356 13574 24366 13626
rect 24366 13574 24412 13626
rect 24116 13572 24172 13574
rect 24196 13572 24252 13574
rect 24276 13572 24332 13574
rect 24356 13572 24412 13574
rect 24116 12538 24172 12540
rect 24196 12538 24252 12540
rect 24276 12538 24332 12540
rect 24356 12538 24412 12540
rect 24116 12486 24162 12538
rect 24162 12486 24172 12538
rect 24196 12486 24226 12538
rect 24226 12486 24238 12538
rect 24238 12486 24252 12538
rect 24276 12486 24290 12538
rect 24290 12486 24302 12538
rect 24302 12486 24332 12538
rect 24356 12486 24366 12538
rect 24366 12486 24412 12538
rect 24116 12484 24172 12486
rect 24196 12484 24252 12486
rect 24276 12484 24332 12486
rect 24356 12484 24412 12486
rect 24858 15036 24860 15056
rect 24860 15036 24912 15056
rect 24912 15036 24914 15056
rect 24858 15000 24914 15036
rect 28354 23160 28410 23216
rect 28354 17040 28410 17096
rect 28354 16360 28410 16416
rect 28354 15000 28410 15056
rect 24858 13368 24914 13424
rect 24116 11450 24172 11452
rect 24196 11450 24252 11452
rect 24276 11450 24332 11452
rect 24356 11450 24412 11452
rect 24116 11398 24162 11450
rect 24162 11398 24172 11450
rect 24196 11398 24226 11450
rect 24226 11398 24238 11450
rect 24238 11398 24252 11450
rect 24276 11398 24290 11450
rect 24290 11398 24302 11450
rect 24302 11398 24332 11450
rect 24356 11398 24366 11450
rect 24366 11398 24412 11450
rect 24116 11396 24172 11398
rect 24196 11396 24252 11398
rect 24276 11396 24332 11398
rect 24356 11396 24412 11398
rect 24116 10362 24172 10364
rect 24196 10362 24252 10364
rect 24276 10362 24332 10364
rect 24356 10362 24412 10364
rect 24116 10310 24162 10362
rect 24162 10310 24172 10362
rect 24196 10310 24226 10362
rect 24226 10310 24238 10362
rect 24238 10310 24252 10362
rect 24276 10310 24290 10362
rect 24290 10310 24302 10362
rect 24302 10310 24332 10362
rect 24356 10310 24366 10362
rect 24366 10310 24412 10362
rect 24116 10308 24172 10310
rect 24196 10308 24252 10310
rect 24276 10308 24332 10310
rect 24356 10308 24412 10310
rect 24116 9274 24172 9276
rect 24196 9274 24252 9276
rect 24276 9274 24332 9276
rect 24356 9274 24412 9276
rect 24116 9222 24162 9274
rect 24162 9222 24172 9274
rect 24196 9222 24226 9274
rect 24226 9222 24238 9274
rect 24238 9222 24252 9274
rect 24276 9222 24290 9274
rect 24290 9222 24302 9274
rect 24302 9222 24332 9274
rect 24356 9222 24366 9274
rect 24366 9222 24412 9274
rect 24116 9220 24172 9222
rect 24196 9220 24252 9222
rect 24276 9220 24332 9222
rect 24356 9220 24412 9222
rect 24116 8186 24172 8188
rect 24196 8186 24252 8188
rect 24276 8186 24332 8188
rect 24356 8186 24412 8188
rect 24116 8134 24162 8186
rect 24162 8134 24172 8186
rect 24196 8134 24226 8186
rect 24226 8134 24238 8186
rect 24238 8134 24252 8186
rect 24276 8134 24290 8186
rect 24290 8134 24302 8186
rect 24302 8134 24332 8186
rect 24356 8134 24366 8186
rect 24366 8134 24412 8186
rect 24116 8132 24172 8134
rect 24196 8132 24252 8134
rect 24276 8132 24332 8134
rect 24356 8132 24412 8134
rect 28262 13640 28318 13696
rect 28354 12280 28410 12336
rect 28262 11600 28318 11656
rect 28262 10240 28318 10296
rect 28354 8916 28356 8936
rect 28356 8916 28408 8936
rect 28408 8916 28410 8936
rect 24116 7098 24172 7100
rect 24196 7098 24252 7100
rect 24276 7098 24332 7100
rect 24356 7098 24412 7100
rect 24116 7046 24162 7098
rect 24162 7046 24172 7098
rect 24196 7046 24226 7098
rect 24226 7046 24238 7098
rect 24238 7046 24252 7098
rect 24276 7046 24290 7098
rect 24290 7046 24302 7098
rect 24302 7046 24332 7098
rect 24356 7046 24366 7098
rect 24366 7046 24412 7098
rect 24116 7044 24172 7046
rect 24196 7044 24252 7046
rect 24276 7044 24332 7046
rect 24356 7044 24412 7046
rect 24116 6010 24172 6012
rect 24196 6010 24252 6012
rect 24276 6010 24332 6012
rect 24356 6010 24412 6012
rect 24116 5958 24162 6010
rect 24162 5958 24172 6010
rect 24196 5958 24226 6010
rect 24226 5958 24238 6010
rect 24238 5958 24252 6010
rect 24276 5958 24290 6010
rect 24290 5958 24302 6010
rect 24302 5958 24332 6010
rect 24356 5958 24366 6010
rect 24366 5958 24412 6010
rect 24116 5956 24172 5958
rect 24196 5956 24252 5958
rect 24276 5956 24332 5958
rect 24356 5956 24412 5958
rect 28354 8880 28410 8916
rect 28354 7520 28410 7576
rect 28354 5480 28410 5536
rect 24116 4922 24172 4924
rect 24196 4922 24252 4924
rect 24276 4922 24332 4924
rect 24356 4922 24412 4924
rect 24116 4870 24162 4922
rect 24162 4870 24172 4922
rect 24196 4870 24226 4922
rect 24226 4870 24238 4922
rect 24238 4870 24252 4922
rect 24276 4870 24290 4922
rect 24290 4870 24302 4922
rect 24302 4870 24332 4922
rect 24356 4870 24366 4922
rect 24366 4870 24412 4922
rect 24116 4868 24172 4870
rect 24196 4868 24252 4870
rect 24276 4868 24332 4870
rect 24356 4868 24412 4870
rect 24116 3834 24172 3836
rect 24196 3834 24252 3836
rect 24276 3834 24332 3836
rect 24356 3834 24412 3836
rect 24116 3782 24162 3834
rect 24162 3782 24172 3834
rect 24196 3782 24226 3834
rect 24226 3782 24238 3834
rect 24238 3782 24252 3834
rect 24276 3782 24290 3834
rect 24290 3782 24302 3834
rect 24302 3782 24332 3834
rect 24356 3782 24366 3834
rect 24366 3782 24412 3834
rect 24116 3780 24172 3782
rect 24196 3780 24252 3782
rect 24276 3780 24332 3782
rect 24356 3780 24412 3782
rect 24116 2746 24172 2748
rect 24196 2746 24252 2748
rect 24276 2746 24332 2748
rect 24356 2746 24412 2748
rect 24116 2694 24162 2746
rect 24162 2694 24172 2746
rect 24196 2694 24226 2746
rect 24226 2694 24238 2746
rect 24238 2694 24252 2746
rect 24276 2694 24290 2746
rect 24290 2694 24302 2746
rect 24302 2694 24332 2746
rect 24356 2694 24366 2746
rect 24366 2694 24412 2746
rect 24116 2692 24172 2694
rect 24196 2692 24252 2694
rect 24276 2692 24332 2694
rect 24356 2692 24412 2694
rect 28354 4120 28410 4176
rect 19484 2202 19540 2204
rect 19564 2202 19620 2204
rect 19644 2202 19700 2204
rect 19724 2202 19780 2204
rect 19484 2150 19530 2202
rect 19530 2150 19540 2202
rect 19564 2150 19594 2202
rect 19594 2150 19606 2202
rect 19606 2150 19620 2202
rect 19644 2150 19658 2202
rect 19658 2150 19670 2202
rect 19670 2150 19700 2202
rect 19724 2150 19734 2202
rect 19734 2150 19780 2202
rect 19484 2148 19540 2150
rect 19564 2148 19620 2150
rect 19644 2148 19700 2150
rect 19724 2148 19780 2150
rect 1674 720 1730 776
rect 28262 720 28318 776
<< metal3 >>
rect 0 29248 800 29368
rect 27521 29338 27587 29341
rect 29200 29338 30000 29368
rect 27521 29336 30000 29338
rect 27521 29280 27526 29336
rect 27582 29280 30000 29336
rect 27521 29278 30000 29280
rect 27521 29275 27587 29278
rect 29200 29248 30000 29278
rect 0 27978 800 28008
rect 1669 27978 1735 27981
rect 0 27976 1735 27978
rect 0 27920 1674 27976
rect 1730 27920 1735 27976
rect 0 27918 1735 27920
rect 0 27888 800 27918
rect 1669 27915 1735 27918
rect 28257 27978 28323 27981
rect 29200 27978 30000 28008
rect 28257 27976 30000 27978
rect 28257 27920 28262 27976
rect 28318 27920 30000 27976
rect 28257 27918 30000 27920
rect 28257 27915 28323 27918
rect 29200 27888 30000 27918
rect 5576 27776 5896 27777
rect 5576 27712 5584 27776
rect 5648 27712 5664 27776
rect 5728 27712 5744 27776
rect 5808 27712 5824 27776
rect 5888 27712 5896 27776
rect 5576 27711 5896 27712
rect 14840 27776 15160 27777
rect 14840 27712 14848 27776
rect 14912 27712 14928 27776
rect 14992 27712 15008 27776
rect 15072 27712 15088 27776
rect 15152 27712 15160 27776
rect 14840 27711 15160 27712
rect 24104 27776 24424 27777
rect 24104 27712 24112 27776
rect 24176 27712 24192 27776
rect 24256 27712 24272 27776
rect 24336 27712 24352 27776
rect 24416 27712 24424 27776
rect 24104 27711 24424 27712
rect 10208 27232 10528 27233
rect 10208 27168 10216 27232
rect 10280 27168 10296 27232
rect 10360 27168 10376 27232
rect 10440 27168 10456 27232
rect 10520 27168 10528 27232
rect 10208 27167 10528 27168
rect 19472 27232 19792 27233
rect 19472 27168 19480 27232
rect 19544 27168 19560 27232
rect 19624 27168 19640 27232
rect 19704 27168 19720 27232
rect 19784 27168 19792 27232
rect 19472 27167 19792 27168
rect 5576 26688 5896 26689
rect 0 26618 800 26648
rect 5576 26624 5584 26688
rect 5648 26624 5664 26688
rect 5728 26624 5744 26688
rect 5808 26624 5824 26688
rect 5888 26624 5896 26688
rect 5576 26623 5896 26624
rect 14840 26688 15160 26689
rect 14840 26624 14848 26688
rect 14912 26624 14928 26688
rect 14992 26624 15008 26688
rect 15072 26624 15088 26688
rect 15152 26624 15160 26688
rect 14840 26623 15160 26624
rect 24104 26688 24424 26689
rect 24104 26624 24112 26688
rect 24176 26624 24192 26688
rect 24256 26624 24272 26688
rect 24336 26624 24352 26688
rect 24416 26624 24424 26688
rect 24104 26623 24424 26624
rect 1393 26618 1459 26621
rect 0 26616 1459 26618
rect 0 26560 1398 26616
rect 1454 26560 1459 26616
rect 0 26558 1459 26560
rect 0 26528 800 26558
rect 1393 26555 1459 26558
rect 28349 26618 28415 26621
rect 29200 26618 30000 26648
rect 28349 26616 30000 26618
rect 28349 26560 28354 26616
rect 28410 26560 30000 26616
rect 28349 26558 30000 26560
rect 28349 26555 28415 26558
rect 29200 26528 30000 26558
rect 10208 26144 10528 26145
rect 10208 26080 10216 26144
rect 10280 26080 10296 26144
rect 10360 26080 10376 26144
rect 10440 26080 10456 26144
rect 10520 26080 10528 26144
rect 10208 26079 10528 26080
rect 19472 26144 19792 26145
rect 19472 26080 19480 26144
rect 19544 26080 19560 26144
rect 19624 26080 19640 26144
rect 19704 26080 19720 26144
rect 19784 26080 19792 26144
rect 19472 26079 19792 26080
rect 0 25938 800 25968
rect 1393 25938 1459 25941
rect 0 25936 1459 25938
rect 0 25880 1398 25936
rect 1454 25880 1459 25936
rect 0 25878 1459 25880
rect 0 25848 800 25878
rect 1393 25875 1459 25878
rect 5576 25600 5896 25601
rect 5576 25536 5584 25600
rect 5648 25536 5664 25600
rect 5728 25536 5744 25600
rect 5808 25536 5824 25600
rect 5888 25536 5896 25600
rect 5576 25535 5896 25536
rect 14840 25600 15160 25601
rect 14840 25536 14848 25600
rect 14912 25536 14928 25600
rect 14992 25536 15008 25600
rect 15072 25536 15088 25600
rect 15152 25536 15160 25600
rect 14840 25535 15160 25536
rect 24104 25600 24424 25601
rect 24104 25536 24112 25600
rect 24176 25536 24192 25600
rect 24256 25536 24272 25600
rect 24336 25536 24352 25600
rect 24416 25536 24424 25600
rect 24104 25535 24424 25536
rect 28349 25258 28415 25261
rect 29200 25258 30000 25288
rect 28349 25256 30000 25258
rect 28349 25200 28354 25256
rect 28410 25200 30000 25256
rect 28349 25198 30000 25200
rect 28349 25195 28415 25198
rect 29200 25168 30000 25198
rect 10208 25056 10528 25057
rect 10208 24992 10216 25056
rect 10280 24992 10296 25056
rect 10360 24992 10376 25056
rect 10440 24992 10456 25056
rect 10520 24992 10528 25056
rect 10208 24991 10528 24992
rect 19472 25056 19792 25057
rect 19472 24992 19480 25056
rect 19544 24992 19560 25056
rect 19624 24992 19640 25056
rect 19704 24992 19720 25056
rect 19784 24992 19792 25056
rect 19472 24991 19792 24992
rect 0 24578 800 24608
rect 1393 24578 1459 24581
rect 0 24576 1459 24578
rect 0 24520 1398 24576
rect 1454 24520 1459 24576
rect 0 24518 1459 24520
rect 0 24488 800 24518
rect 1393 24515 1459 24518
rect 5576 24512 5896 24513
rect 5576 24448 5584 24512
rect 5648 24448 5664 24512
rect 5728 24448 5744 24512
rect 5808 24448 5824 24512
rect 5888 24448 5896 24512
rect 5576 24447 5896 24448
rect 14840 24512 15160 24513
rect 14840 24448 14848 24512
rect 14912 24448 14928 24512
rect 14992 24448 15008 24512
rect 15072 24448 15088 24512
rect 15152 24448 15160 24512
rect 14840 24447 15160 24448
rect 24104 24512 24424 24513
rect 24104 24448 24112 24512
rect 24176 24448 24192 24512
rect 24256 24448 24272 24512
rect 24336 24448 24352 24512
rect 24416 24448 24424 24512
rect 29200 24488 30000 24608
rect 24104 24447 24424 24448
rect 10208 23968 10528 23969
rect 10208 23904 10216 23968
rect 10280 23904 10296 23968
rect 10360 23904 10376 23968
rect 10440 23904 10456 23968
rect 10520 23904 10528 23968
rect 10208 23903 10528 23904
rect 19472 23968 19792 23969
rect 19472 23904 19480 23968
rect 19544 23904 19560 23968
rect 19624 23904 19640 23968
rect 19704 23904 19720 23968
rect 19784 23904 19792 23968
rect 19472 23903 19792 23904
rect 5576 23424 5896 23425
rect 5576 23360 5584 23424
rect 5648 23360 5664 23424
rect 5728 23360 5744 23424
rect 5808 23360 5824 23424
rect 5888 23360 5896 23424
rect 5576 23359 5896 23360
rect 14840 23424 15160 23425
rect 14840 23360 14848 23424
rect 14912 23360 14928 23424
rect 14992 23360 15008 23424
rect 15072 23360 15088 23424
rect 15152 23360 15160 23424
rect 14840 23359 15160 23360
rect 24104 23424 24424 23425
rect 24104 23360 24112 23424
rect 24176 23360 24192 23424
rect 24256 23360 24272 23424
rect 24336 23360 24352 23424
rect 24416 23360 24424 23424
rect 24104 23359 24424 23360
rect 0 23218 800 23248
rect 1393 23218 1459 23221
rect 0 23216 1459 23218
rect 0 23160 1398 23216
rect 1454 23160 1459 23216
rect 0 23158 1459 23160
rect 0 23128 800 23158
rect 1393 23155 1459 23158
rect 28349 23218 28415 23221
rect 29200 23218 30000 23248
rect 28349 23216 30000 23218
rect 28349 23160 28354 23216
rect 28410 23160 30000 23216
rect 28349 23158 30000 23160
rect 28349 23155 28415 23158
rect 29200 23128 30000 23158
rect 10208 22880 10528 22881
rect 10208 22816 10216 22880
rect 10280 22816 10296 22880
rect 10360 22816 10376 22880
rect 10440 22816 10456 22880
rect 10520 22816 10528 22880
rect 10208 22815 10528 22816
rect 19472 22880 19792 22881
rect 19472 22816 19480 22880
rect 19544 22816 19560 22880
rect 19624 22816 19640 22880
rect 19704 22816 19720 22880
rect 19784 22816 19792 22880
rect 19472 22815 19792 22816
rect 5576 22336 5896 22337
rect 5576 22272 5584 22336
rect 5648 22272 5664 22336
rect 5728 22272 5744 22336
rect 5808 22272 5824 22336
rect 5888 22272 5896 22336
rect 5576 22271 5896 22272
rect 14840 22336 15160 22337
rect 14840 22272 14848 22336
rect 14912 22272 14928 22336
rect 14992 22272 15008 22336
rect 15072 22272 15088 22336
rect 15152 22272 15160 22336
rect 14840 22271 15160 22272
rect 24104 22336 24424 22337
rect 24104 22272 24112 22336
rect 24176 22272 24192 22336
rect 24256 22272 24272 22336
rect 24336 22272 24352 22336
rect 24416 22272 24424 22336
rect 24104 22271 24424 22272
rect 0 21768 800 21888
rect 10208 21792 10528 21793
rect 10208 21728 10216 21792
rect 10280 21728 10296 21792
rect 10360 21728 10376 21792
rect 10440 21728 10456 21792
rect 10520 21728 10528 21792
rect 10208 21727 10528 21728
rect 19472 21792 19792 21793
rect 19472 21728 19480 21792
rect 19544 21728 19560 21792
rect 19624 21728 19640 21792
rect 19704 21728 19720 21792
rect 19784 21728 19792 21792
rect 29200 21768 30000 21888
rect 19472 21727 19792 21728
rect 17217 21314 17283 21317
rect 17534 21314 17540 21316
rect 17217 21312 17540 21314
rect 17217 21256 17222 21312
rect 17278 21256 17540 21312
rect 17217 21254 17540 21256
rect 17217 21251 17283 21254
rect 17534 21252 17540 21254
rect 17604 21314 17610 21316
rect 19333 21314 19399 21317
rect 17604 21312 19399 21314
rect 17604 21256 19338 21312
rect 19394 21256 19399 21312
rect 17604 21254 19399 21256
rect 17604 21252 17610 21254
rect 19333 21251 19399 21254
rect 5576 21248 5896 21249
rect 0 21178 800 21208
rect 5576 21184 5584 21248
rect 5648 21184 5664 21248
rect 5728 21184 5744 21248
rect 5808 21184 5824 21248
rect 5888 21184 5896 21248
rect 5576 21183 5896 21184
rect 14840 21248 15160 21249
rect 14840 21184 14848 21248
rect 14912 21184 14928 21248
rect 14992 21184 15008 21248
rect 15072 21184 15088 21248
rect 15152 21184 15160 21248
rect 14840 21183 15160 21184
rect 24104 21248 24424 21249
rect 24104 21184 24112 21248
rect 24176 21184 24192 21248
rect 24256 21184 24272 21248
rect 24336 21184 24352 21248
rect 24416 21184 24424 21248
rect 24104 21183 24424 21184
rect 1393 21178 1459 21181
rect 0 21176 1459 21178
rect 0 21120 1398 21176
rect 1454 21120 1459 21176
rect 0 21118 1459 21120
rect 0 21088 800 21118
rect 1393 21115 1459 21118
rect 29200 21088 30000 21208
rect 10208 20704 10528 20705
rect 10208 20640 10216 20704
rect 10280 20640 10296 20704
rect 10360 20640 10376 20704
rect 10440 20640 10456 20704
rect 10520 20640 10528 20704
rect 10208 20639 10528 20640
rect 19472 20704 19792 20705
rect 19472 20640 19480 20704
rect 19544 20640 19560 20704
rect 19624 20640 19640 20704
rect 19704 20640 19720 20704
rect 19784 20640 19792 20704
rect 19472 20639 19792 20640
rect 5576 20160 5896 20161
rect 5576 20096 5584 20160
rect 5648 20096 5664 20160
rect 5728 20096 5744 20160
rect 5808 20096 5824 20160
rect 5888 20096 5896 20160
rect 5576 20095 5896 20096
rect 14840 20160 15160 20161
rect 14840 20096 14848 20160
rect 14912 20096 14928 20160
rect 14992 20096 15008 20160
rect 15072 20096 15088 20160
rect 15152 20096 15160 20160
rect 14840 20095 15160 20096
rect 24104 20160 24424 20161
rect 24104 20096 24112 20160
rect 24176 20096 24192 20160
rect 24256 20096 24272 20160
rect 24336 20096 24352 20160
rect 24416 20096 24424 20160
rect 24104 20095 24424 20096
rect 0 19818 800 19848
rect 1393 19818 1459 19821
rect 0 19816 1459 19818
rect 0 19760 1398 19816
rect 1454 19760 1459 19816
rect 0 19758 1459 19760
rect 0 19728 800 19758
rect 1393 19755 1459 19758
rect 29200 19728 30000 19848
rect 21081 19684 21147 19685
rect 21030 19620 21036 19684
rect 21100 19682 21147 19684
rect 21100 19680 21192 19682
rect 21142 19624 21192 19680
rect 21100 19622 21192 19624
rect 21100 19620 21147 19622
rect 21081 19619 21147 19620
rect 10208 19616 10528 19617
rect 10208 19552 10216 19616
rect 10280 19552 10296 19616
rect 10360 19552 10376 19616
rect 10440 19552 10456 19616
rect 10520 19552 10528 19616
rect 10208 19551 10528 19552
rect 19472 19616 19792 19617
rect 19472 19552 19480 19616
rect 19544 19552 19560 19616
rect 19624 19552 19640 19616
rect 19704 19552 19720 19616
rect 19784 19552 19792 19616
rect 19472 19551 19792 19552
rect 5576 19072 5896 19073
rect 5576 19008 5584 19072
rect 5648 19008 5664 19072
rect 5728 19008 5744 19072
rect 5808 19008 5824 19072
rect 5888 19008 5896 19072
rect 5576 19007 5896 19008
rect 14840 19072 15160 19073
rect 14840 19008 14848 19072
rect 14912 19008 14928 19072
rect 14992 19008 15008 19072
rect 15072 19008 15088 19072
rect 15152 19008 15160 19072
rect 14840 19007 15160 19008
rect 24104 19072 24424 19073
rect 24104 19008 24112 19072
rect 24176 19008 24192 19072
rect 24256 19008 24272 19072
rect 24336 19008 24352 19072
rect 24416 19008 24424 19072
rect 24104 19007 24424 19008
rect 10208 18528 10528 18529
rect 0 18458 800 18488
rect 10208 18464 10216 18528
rect 10280 18464 10296 18528
rect 10360 18464 10376 18528
rect 10440 18464 10456 18528
rect 10520 18464 10528 18528
rect 10208 18463 10528 18464
rect 19472 18528 19792 18529
rect 19472 18464 19480 18528
rect 19544 18464 19560 18528
rect 19624 18464 19640 18528
rect 19704 18464 19720 18528
rect 19784 18464 19792 18528
rect 19472 18463 19792 18464
rect 1393 18458 1459 18461
rect 0 18456 1459 18458
rect 0 18400 1398 18456
rect 1454 18400 1459 18456
rect 0 18398 1459 18400
rect 0 18368 800 18398
rect 1393 18395 1459 18398
rect 29200 18368 30000 18488
rect 5576 17984 5896 17985
rect 5576 17920 5584 17984
rect 5648 17920 5664 17984
rect 5728 17920 5744 17984
rect 5808 17920 5824 17984
rect 5888 17920 5896 17984
rect 5576 17919 5896 17920
rect 14840 17984 15160 17985
rect 14840 17920 14848 17984
rect 14912 17920 14928 17984
rect 14992 17920 15008 17984
rect 15072 17920 15088 17984
rect 15152 17920 15160 17984
rect 14840 17919 15160 17920
rect 24104 17984 24424 17985
rect 24104 17920 24112 17984
rect 24176 17920 24192 17984
rect 24256 17920 24272 17984
rect 24336 17920 24352 17984
rect 24416 17920 24424 17984
rect 24104 17919 24424 17920
rect 16481 17642 16547 17645
rect 22093 17642 22159 17645
rect 16481 17640 22159 17642
rect 16481 17584 16486 17640
rect 16542 17584 22098 17640
rect 22154 17584 22159 17640
rect 16481 17582 22159 17584
rect 16481 17579 16547 17582
rect 22093 17579 22159 17582
rect 10208 17440 10528 17441
rect 10208 17376 10216 17440
rect 10280 17376 10296 17440
rect 10360 17376 10376 17440
rect 10440 17376 10456 17440
rect 10520 17376 10528 17440
rect 10208 17375 10528 17376
rect 19472 17440 19792 17441
rect 19472 17376 19480 17440
rect 19544 17376 19560 17440
rect 19624 17376 19640 17440
rect 19704 17376 19720 17440
rect 19784 17376 19792 17440
rect 19472 17375 19792 17376
rect 1761 17234 1827 17237
rect 18321 17234 18387 17237
rect 1761 17232 18387 17234
rect 1761 17176 1766 17232
rect 1822 17176 18326 17232
rect 18382 17176 18387 17232
rect 1761 17174 18387 17176
rect 1761 17171 1827 17174
rect 18321 17171 18387 17174
rect 0 17098 800 17128
rect 1393 17098 1459 17101
rect 0 17096 1459 17098
rect 0 17040 1398 17096
rect 1454 17040 1459 17096
rect 0 17038 1459 17040
rect 0 17008 800 17038
rect 1393 17035 1459 17038
rect 12709 17098 12775 17101
rect 14457 17098 14523 17101
rect 12709 17096 14523 17098
rect 12709 17040 12714 17096
rect 12770 17040 14462 17096
rect 14518 17040 14523 17096
rect 12709 17038 14523 17040
rect 12709 17035 12775 17038
rect 14457 17035 14523 17038
rect 28349 17098 28415 17101
rect 29200 17098 30000 17128
rect 28349 17096 30000 17098
rect 28349 17040 28354 17096
rect 28410 17040 30000 17096
rect 28349 17038 30000 17040
rect 28349 17035 28415 17038
rect 29200 17008 30000 17038
rect 14365 16962 14431 16965
rect 14365 16960 14474 16962
rect 14365 16904 14370 16960
rect 14426 16904 14474 16960
rect 14365 16899 14474 16904
rect 5576 16896 5896 16897
rect 5576 16832 5584 16896
rect 5648 16832 5664 16896
rect 5728 16832 5744 16896
rect 5808 16832 5824 16896
rect 5888 16832 5896 16896
rect 5576 16831 5896 16832
rect 14414 16693 14474 16899
rect 14840 16896 15160 16897
rect 14840 16832 14848 16896
rect 14912 16832 14928 16896
rect 14992 16832 15008 16896
rect 15072 16832 15088 16896
rect 15152 16832 15160 16896
rect 14840 16831 15160 16832
rect 24104 16896 24424 16897
rect 24104 16832 24112 16896
rect 24176 16832 24192 16896
rect 24256 16832 24272 16896
rect 24336 16832 24352 16896
rect 24416 16832 24424 16896
rect 24104 16831 24424 16832
rect 13813 16692 13879 16693
rect 13813 16688 13860 16692
rect 13924 16690 13930 16692
rect 14089 16690 14155 16693
rect 14222 16690 14228 16692
rect 13813 16632 13818 16688
rect 13813 16628 13860 16632
rect 13924 16630 13970 16690
rect 14089 16688 14228 16690
rect 14089 16632 14094 16688
rect 14150 16632 14228 16688
rect 14089 16630 14228 16632
rect 13924 16628 13930 16630
rect 13813 16627 13879 16628
rect 14089 16627 14155 16630
rect 14222 16628 14228 16630
rect 14292 16628 14298 16692
rect 14414 16688 14523 16693
rect 14414 16632 14462 16688
rect 14518 16632 14523 16688
rect 14414 16630 14523 16632
rect 14457 16627 14523 16630
rect 13353 16554 13419 16557
rect 15377 16554 15443 16557
rect 13353 16552 15443 16554
rect 13353 16496 13358 16552
rect 13414 16496 15382 16552
rect 15438 16496 15443 16552
rect 13353 16494 15443 16496
rect 13353 16491 13419 16494
rect 15377 16491 15443 16494
rect 0 16418 800 16448
rect 1485 16418 1551 16421
rect 0 16416 1551 16418
rect 0 16360 1490 16416
rect 1546 16360 1551 16416
rect 0 16358 1551 16360
rect 0 16328 800 16358
rect 1485 16355 1551 16358
rect 12893 16418 12959 16421
rect 13997 16418 14063 16421
rect 12893 16416 14063 16418
rect 12893 16360 12898 16416
rect 12954 16360 14002 16416
rect 14058 16360 14063 16416
rect 12893 16358 14063 16360
rect 12893 16355 12959 16358
rect 13997 16355 14063 16358
rect 14181 16418 14247 16421
rect 15193 16418 15259 16421
rect 14181 16416 15259 16418
rect 14181 16360 14186 16416
rect 14242 16360 15198 16416
rect 15254 16360 15259 16416
rect 14181 16358 15259 16360
rect 14181 16355 14247 16358
rect 15193 16355 15259 16358
rect 28349 16418 28415 16421
rect 29200 16418 30000 16448
rect 28349 16416 30000 16418
rect 28349 16360 28354 16416
rect 28410 16360 30000 16416
rect 28349 16358 30000 16360
rect 28349 16355 28415 16358
rect 10208 16352 10528 16353
rect 10208 16288 10216 16352
rect 10280 16288 10296 16352
rect 10360 16288 10376 16352
rect 10440 16288 10456 16352
rect 10520 16288 10528 16352
rect 10208 16287 10528 16288
rect 19472 16352 19792 16353
rect 19472 16288 19480 16352
rect 19544 16288 19560 16352
rect 19624 16288 19640 16352
rect 19704 16288 19720 16352
rect 19784 16288 19792 16352
rect 29200 16328 30000 16358
rect 19472 16287 19792 16288
rect 13537 16282 13603 16285
rect 19333 16282 19399 16285
rect 13537 16280 19399 16282
rect 13537 16224 13542 16280
rect 13598 16224 19338 16280
rect 19394 16224 19399 16280
rect 13537 16222 19399 16224
rect 13537 16219 13603 16222
rect 19333 16219 19399 16222
rect 14549 16146 14615 16149
rect 20989 16146 21055 16149
rect 14549 16144 21055 16146
rect 14549 16088 14554 16144
rect 14610 16088 20994 16144
rect 21050 16088 21055 16144
rect 14549 16086 21055 16088
rect 14549 16083 14615 16086
rect 20989 16083 21055 16086
rect 15377 16010 15443 16013
rect 22093 16010 22159 16013
rect 15377 16008 22159 16010
rect 15377 15952 15382 16008
rect 15438 15952 22098 16008
rect 22154 15952 22159 16008
rect 15377 15950 22159 15952
rect 15377 15947 15443 15950
rect 22093 15947 22159 15950
rect 5576 15808 5896 15809
rect 5576 15744 5584 15808
rect 5648 15744 5664 15808
rect 5728 15744 5744 15808
rect 5808 15744 5824 15808
rect 5888 15744 5896 15808
rect 5576 15743 5896 15744
rect 14840 15808 15160 15809
rect 14840 15744 14848 15808
rect 14912 15744 14928 15808
rect 14992 15744 15008 15808
rect 15072 15744 15088 15808
rect 15152 15744 15160 15808
rect 14840 15743 15160 15744
rect 24104 15808 24424 15809
rect 24104 15744 24112 15808
rect 24176 15744 24192 15808
rect 24256 15744 24272 15808
rect 24336 15744 24352 15808
rect 24416 15744 24424 15808
rect 24104 15743 24424 15744
rect 13997 15602 14063 15605
rect 15377 15602 15443 15605
rect 13997 15600 15443 15602
rect 13997 15544 14002 15600
rect 14058 15544 15382 15600
rect 15438 15544 15443 15600
rect 13997 15542 15443 15544
rect 13997 15539 14063 15542
rect 15377 15539 15443 15542
rect 10961 15466 11027 15469
rect 12985 15466 13051 15469
rect 17125 15466 17191 15469
rect 21030 15466 21036 15468
rect 10961 15464 21036 15466
rect 10961 15408 10966 15464
rect 11022 15408 12990 15464
rect 13046 15408 17130 15464
rect 17186 15408 21036 15464
rect 10961 15406 21036 15408
rect 10961 15403 11027 15406
rect 12985 15403 13051 15406
rect 17125 15403 17191 15406
rect 21030 15404 21036 15406
rect 21100 15466 21106 15468
rect 22001 15466 22067 15469
rect 21100 15464 22067 15466
rect 21100 15408 22006 15464
rect 22062 15408 22067 15464
rect 21100 15406 22067 15408
rect 21100 15404 21106 15406
rect 22001 15403 22067 15406
rect 10208 15264 10528 15265
rect 10208 15200 10216 15264
rect 10280 15200 10296 15264
rect 10360 15200 10376 15264
rect 10440 15200 10456 15264
rect 10520 15200 10528 15264
rect 10208 15199 10528 15200
rect 19472 15264 19792 15265
rect 19472 15200 19480 15264
rect 19544 15200 19560 15264
rect 19624 15200 19640 15264
rect 19704 15200 19720 15264
rect 19784 15200 19792 15264
rect 19472 15199 19792 15200
rect 20437 15194 20503 15197
rect 23841 15194 23907 15197
rect 20437 15192 23907 15194
rect 20437 15136 20442 15192
rect 20498 15136 23846 15192
rect 23902 15136 23907 15192
rect 20437 15134 23907 15136
rect 20437 15131 20503 15134
rect 23841 15131 23907 15134
rect 0 14968 800 15088
rect 16205 15058 16271 15061
rect 16941 15058 17007 15061
rect 17677 15058 17743 15061
rect 16205 15056 17743 15058
rect 16205 15000 16210 15056
rect 16266 15000 16946 15056
rect 17002 15000 17682 15056
rect 17738 15000 17743 15056
rect 16205 14998 17743 15000
rect 16205 14995 16271 14998
rect 16941 14995 17007 14998
rect 17677 14995 17743 14998
rect 17861 15058 17927 15061
rect 19793 15058 19859 15061
rect 17861 15056 19859 15058
rect 17861 15000 17866 15056
rect 17922 15000 19798 15056
rect 19854 15000 19859 15056
rect 17861 14998 19859 15000
rect 17861 14995 17927 14998
rect 19793 14995 19859 14998
rect 20713 15058 20779 15061
rect 24853 15058 24919 15061
rect 20713 15056 24919 15058
rect 20713 15000 20718 15056
rect 20774 15000 24858 15056
rect 24914 15000 24919 15056
rect 20713 14998 24919 15000
rect 20713 14995 20779 14998
rect 24853 14995 24919 14998
rect 28349 15058 28415 15061
rect 29200 15058 30000 15088
rect 28349 15056 30000 15058
rect 28349 15000 28354 15056
rect 28410 15000 30000 15056
rect 28349 14998 30000 15000
rect 28349 14995 28415 14998
rect 29200 14968 30000 14998
rect 14273 14922 14339 14925
rect 14457 14922 14523 14925
rect 23473 14922 23539 14925
rect 14273 14920 23539 14922
rect 14273 14864 14278 14920
rect 14334 14864 14462 14920
rect 14518 14864 23478 14920
rect 23534 14864 23539 14920
rect 14273 14862 23539 14864
rect 14273 14859 14339 14862
rect 14457 14859 14523 14862
rect 23473 14859 23539 14862
rect 5576 14720 5896 14721
rect 5576 14656 5584 14720
rect 5648 14656 5664 14720
rect 5728 14656 5744 14720
rect 5808 14656 5824 14720
rect 5888 14656 5896 14720
rect 5576 14655 5896 14656
rect 14840 14720 15160 14721
rect 14840 14656 14848 14720
rect 14912 14656 14928 14720
rect 14992 14656 15008 14720
rect 15072 14656 15088 14720
rect 15152 14656 15160 14720
rect 14840 14655 15160 14656
rect 24104 14720 24424 14721
rect 24104 14656 24112 14720
rect 24176 14656 24192 14720
rect 24256 14656 24272 14720
rect 24336 14656 24352 14720
rect 24416 14656 24424 14720
rect 24104 14655 24424 14656
rect 13261 14514 13327 14517
rect 15193 14514 15259 14517
rect 15326 14514 15332 14516
rect 13261 14512 15332 14514
rect 13261 14456 13266 14512
rect 13322 14456 15198 14512
rect 15254 14456 15332 14512
rect 13261 14454 15332 14456
rect 13261 14451 13327 14454
rect 15193 14451 15259 14454
rect 15326 14452 15332 14454
rect 15396 14452 15402 14516
rect 13169 14378 13235 14381
rect 17033 14378 17099 14381
rect 13169 14376 17099 14378
rect 13169 14320 13174 14376
rect 13230 14320 17038 14376
rect 17094 14320 17099 14376
rect 13169 14318 17099 14320
rect 13169 14315 13235 14318
rect 17033 14315 17099 14318
rect 10208 14176 10528 14177
rect 10208 14112 10216 14176
rect 10280 14112 10296 14176
rect 10360 14112 10376 14176
rect 10440 14112 10456 14176
rect 10520 14112 10528 14176
rect 10208 14111 10528 14112
rect 19472 14176 19792 14177
rect 19472 14112 19480 14176
rect 19544 14112 19560 14176
rect 19624 14112 19640 14176
rect 19704 14112 19720 14176
rect 19784 14112 19792 14176
rect 19472 14111 19792 14112
rect 0 13698 800 13728
rect 1393 13698 1459 13701
rect 0 13696 1459 13698
rect 0 13640 1398 13696
rect 1454 13640 1459 13696
rect 0 13638 1459 13640
rect 0 13608 800 13638
rect 1393 13635 1459 13638
rect 9489 13698 9555 13701
rect 13169 13698 13235 13701
rect 9489 13696 13235 13698
rect 9489 13640 9494 13696
rect 9550 13640 13174 13696
rect 13230 13640 13235 13696
rect 9489 13638 13235 13640
rect 9489 13635 9555 13638
rect 13169 13635 13235 13638
rect 28257 13698 28323 13701
rect 29200 13698 30000 13728
rect 28257 13696 30000 13698
rect 28257 13640 28262 13696
rect 28318 13640 30000 13696
rect 28257 13638 30000 13640
rect 28257 13635 28323 13638
rect 5576 13632 5896 13633
rect 5576 13568 5584 13632
rect 5648 13568 5664 13632
rect 5728 13568 5744 13632
rect 5808 13568 5824 13632
rect 5888 13568 5896 13632
rect 5576 13567 5896 13568
rect 14840 13632 15160 13633
rect 14840 13568 14848 13632
rect 14912 13568 14928 13632
rect 14992 13568 15008 13632
rect 15072 13568 15088 13632
rect 15152 13568 15160 13632
rect 14840 13567 15160 13568
rect 24104 13632 24424 13633
rect 24104 13568 24112 13632
rect 24176 13568 24192 13632
rect 24256 13568 24272 13632
rect 24336 13568 24352 13632
rect 24416 13568 24424 13632
rect 29200 13608 30000 13638
rect 24104 13567 24424 13568
rect 17585 13426 17651 13429
rect 24853 13426 24919 13429
rect 17585 13424 24919 13426
rect 17585 13368 17590 13424
rect 17646 13368 24858 13424
rect 24914 13368 24919 13424
rect 17585 13366 24919 13368
rect 17585 13363 17651 13366
rect 24853 13363 24919 13366
rect 15326 13228 15332 13292
rect 15396 13290 15402 13292
rect 22461 13290 22527 13293
rect 15396 13288 22527 13290
rect 15396 13232 22466 13288
rect 22522 13232 22527 13288
rect 15396 13230 22527 13232
rect 15396 13228 15402 13230
rect 22461 13227 22527 13230
rect 10208 13088 10528 13089
rect 0 12928 800 13048
rect 10208 13024 10216 13088
rect 10280 13024 10296 13088
rect 10360 13024 10376 13088
rect 10440 13024 10456 13088
rect 10520 13024 10528 13088
rect 10208 13023 10528 13024
rect 19472 13088 19792 13089
rect 19472 13024 19480 13088
rect 19544 13024 19560 13088
rect 19624 13024 19640 13088
rect 19704 13024 19720 13088
rect 19784 13024 19792 13088
rect 19472 13023 19792 13024
rect 5576 12544 5896 12545
rect 5576 12480 5584 12544
rect 5648 12480 5664 12544
rect 5728 12480 5744 12544
rect 5808 12480 5824 12544
rect 5888 12480 5896 12544
rect 5576 12479 5896 12480
rect 14840 12544 15160 12545
rect 14840 12480 14848 12544
rect 14912 12480 14928 12544
rect 14992 12480 15008 12544
rect 15072 12480 15088 12544
rect 15152 12480 15160 12544
rect 14840 12479 15160 12480
rect 24104 12544 24424 12545
rect 24104 12480 24112 12544
rect 24176 12480 24192 12544
rect 24256 12480 24272 12544
rect 24336 12480 24352 12544
rect 24416 12480 24424 12544
rect 24104 12479 24424 12480
rect 14733 12338 14799 12341
rect 20805 12338 20871 12341
rect 14733 12336 20871 12338
rect 14733 12280 14738 12336
rect 14794 12280 20810 12336
rect 20866 12280 20871 12336
rect 14733 12278 20871 12280
rect 14733 12275 14799 12278
rect 20805 12275 20871 12278
rect 28349 12338 28415 12341
rect 29200 12338 30000 12368
rect 28349 12336 30000 12338
rect 28349 12280 28354 12336
rect 28410 12280 30000 12336
rect 28349 12278 30000 12280
rect 28349 12275 28415 12278
rect 29200 12248 30000 12278
rect 13813 12202 13879 12205
rect 18229 12202 18295 12205
rect 22553 12202 22619 12205
rect 13813 12200 18295 12202
rect 13813 12144 13818 12200
rect 13874 12144 18234 12200
rect 18290 12144 18295 12200
rect 13813 12142 18295 12144
rect 13813 12139 13879 12142
rect 18229 12139 18295 12142
rect 19290 12200 22619 12202
rect 19290 12144 22558 12200
rect 22614 12144 22619 12200
rect 19290 12142 22619 12144
rect 17493 12068 17559 12069
rect 17493 12064 17540 12068
rect 17604 12066 17610 12068
rect 17493 12008 17498 12064
rect 17493 12004 17540 12008
rect 17604 12006 17650 12066
rect 17604 12004 17610 12006
rect 17493 12003 17559 12004
rect 10208 12000 10528 12001
rect 10208 11936 10216 12000
rect 10280 11936 10296 12000
rect 10360 11936 10376 12000
rect 10440 11936 10456 12000
rect 10520 11936 10528 12000
rect 10208 11935 10528 11936
rect 15193 11930 15259 11933
rect 19290 11930 19350 12142
rect 22553 12139 22619 12142
rect 19472 12000 19792 12001
rect 19472 11936 19480 12000
rect 19544 11936 19560 12000
rect 19624 11936 19640 12000
rect 19704 11936 19720 12000
rect 19784 11936 19792 12000
rect 19472 11935 19792 11936
rect 15193 11928 19350 11930
rect 15193 11872 15198 11928
rect 15254 11872 19350 11928
rect 15193 11870 19350 11872
rect 15193 11867 15259 11870
rect 10225 11794 10291 11797
rect 10961 11794 11027 11797
rect 10225 11792 11027 11794
rect 10225 11736 10230 11792
rect 10286 11736 10966 11792
rect 11022 11736 11027 11792
rect 10225 11734 11027 11736
rect 10225 11731 10291 11734
rect 10961 11731 11027 11734
rect 0 11568 800 11688
rect 28257 11658 28323 11661
rect 29200 11658 30000 11688
rect 28257 11656 30000 11658
rect 28257 11600 28262 11656
rect 28318 11600 30000 11656
rect 28257 11598 30000 11600
rect 28257 11595 28323 11598
rect 29200 11568 30000 11598
rect 5576 11456 5896 11457
rect 5576 11392 5584 11456
rect 5648 11392 5664 11456
rect 5728 11392 5744 11456
rect 5808 11392 5824 11456
rect 5888 11392 5896 11456
rect 5576 11391 5896 11392
rect 14840 11456 15160 11457
rect 14840 11392 14848 11456
rect 14912 11392 14928 11456
rect 14992 11392 15008 11456
rect 15072 11392 15088 11456
rect 15152 11392 15160 11456
rect 14840 11391 15160 11392
rect 24104 11456 24424 11457
rect 24104 11392 24112 11456
rect 24176 11392 24192 11456
rect 24256 11392 24272 11456
rect 24336 11392 24352 11456
rect 24416 11392 24424 11456
rect 24104 11391 24424 11392
rect 10317 11250 10383 11253
rect 15009 11250 15075 11253
rect 10317 11248 15075 11250
rect 10317 11192 10322 11248
rect 10378 11192 15014 11248
rect 15070 11192 15075 11248
rect 10317 11190 15075 11192
rect 10317 11187 10383 11190
rect 15009 11187 15075 11190
rect 11145 11116 11211 11117
rect 11094 11114 11100 11116
rect 11054 11054 11100 11114
rect 11164 11112 11211 11116
rect 11206 11056 11211 11112
rect 11094 11052 11100 11054
rect 11164 11052 11211 11056
rect 11145 11051 11211 11052
rect 10208 10912 10528 10913
rect 10208 10848 10216 10912
rect 10280 10848 10296 10912
rect 10360 10848 10376 10912
rect 10440 10848 10456 10912
rect 10520 10848 10528 10912
rect 10208 10847 10528 10848
rect 19472 10912 19792 10913
rect 19472 10848 19480 10912
rect 19544 10848 19560 10912
rect 19624 10848 19640 10912
rect 19704 10848 19720 10912
rect 19784 10848 19792 10912
rect 19472 10847 19792 10848
rect 5576 10368 5896 10369
rect 0 10298 800 10328
rect 5576 10304 5584 10368
rect 5648 10304 5664 10368
rect 5728 10304 5744 10368
rect 5808 10304 5824 10368
rect 5888 10304 5896 10368
rect 5576 10303 5896 10304
rect 14840 10368 15160 10369
rect 14840 10304 14848 10368
rect 14912 10304 14928 10368
rect 14992 10304 15008 10368
rect 15072 10304 15088 10368
rect 15152 10304 15160 10368
rect 14840 10303 15160 10304
rect 24104 10368 24424 10369
rect 24104 10304 24112 10368
rect 24176 10304 24192 10368
rect 24256 10304 24272 10368
rect 24336 10304 24352 10368
rect 24416 10304 24424 10368
rect 24104 10303 24424 10304
rect 1393 10298 1459 10301
rect 0 10296 1459 10298
rect 0 10240 1398 10296
rect 1454 10240 1459 10296
rect 0 10238 1459 10240
rect 0 10208 800 10238
rect 1393 10235 1459 10238
rect 28257 10298 28323 10301
rect 29200 10298 30000 10328
rect 28257 10296 30000 10298
rect 28257 10240 28262 10296
rect 28318 10240 30000 10296
rect 28257 10238 30000 10240
rect 28257 10235 28323 10238
rect 29200 10208 30000 10238
rect 10208 9824 10528 9825
rect 10208 9760 10216 9824
rect 10280 9760 10296 9824
rect 10360 9760 10376 9824
rect 10440 9760 10456 9824
rect 10520 9760 10528 9824
rect 10208 9759 10528 9760
rect 19472 9824 19792 9825
rect 19472 9760 19480 9824
rect 19544 9760 19560 9824
rect 19624 9760 19640 9824
rect 19704 9760 19720 9824
rect 19784 9760 19792 9824
rect 19472 9759 19792 9760
rect 7465 9618 7531 9621
rect 9121 9618 9187 9621
rect 7465 9616 9187 9618
rect 7465 9560 7470 9616
rect 7526 9560 9126 9616
rect 9182 9560 9187 9616
rect 7465 9558 9187 9560
rect 7465 9555 7531 9558
rect 9121 9555 9187 9558
rect 5576 9280 5896 9281
rect 5576 9216 5584 9280
rect 5648 9216 5664 9280
rect 5728 9216 5744 9280
rect 5808 9216 5824 9280
rect 5888 9216 5896 9280
rect 5576 9215 5896 9216
rect 14840 9280 15160 9281
rect 14840 9216 14848 9280
rect 14912 9216 14928 9280
rect 14992 9216 15008 9280
rect 15072 9216 15088 9280
rect 15152 9216 15160 9280
rect 14840 9215 15160 9216
rect 24104 9280 24424 9281
rect 24104 9216 24112 9280
rect 24176 9216 24192 9280
rect 24256 9216 24272 9280
rect 24336 9216 24352 9280
rect 24416 9216 24424 9280
rect 24104 9215 24424 9216
rect 0 8938 800 8968
rect 1669 8938 1735 8941
rect 0 8936 1735 8938
rect 0 8880 1674 8936
rect 1730 8880 1735 8936
rect 0 8878 1735 8880
rect 0 8848 800 8878
rect 1669 8875 1735 8878
rect 1853 8938 1919 8941
rect 16113 8938 16179 8941
rect 1853 8936 16179 8938
rect 1853 8880 1858 8936
rect 1914 8880 16118 8936
rect 16174 8880 16179 8936
rect 1853 8878 16179 8880
rect 1853 8875 1919 8878
rect 16113 8875 16179 8878
rect 28349 8938 28415 8941
rect 29200 8938 30000 8968
rect 28349 8936 30000 8938
rect 28349 8880 28354 8936
rect 28410 8880 30000 8936
rect 28349 8878 30000 8880
rect 28349 8875 28415 8878
rect 29200 8848 30000 8878
rect 10208 8736 10528 8737
rect 10208 8672 10216 8736
rect 10280 8672 10296 8736
rect 10360 8672 10376 8736
rect 10440 8672 10456 8736
rect 10520 8672 10528 8736
rect 10208 8671 10528 8672
rect 19472 8736 19792 8737
rect 19472 8672 19480 8736
rect 19544 8672 19560 8736
rect 19624 8672 19640 8736
rect 19704 8672 19720 8736
rect 19784 8672 19792 8736
rect 19472 8671 19792 8672
rect 9673 8530 9739 8533
rect 12341 8530 12407 8533
rect 9673 8528 12407 8530
rect 9673 8472 9678 8528
rect 9734 8472 12346 8528
rect 12402 8472 12407 8528
rect 9673 8470 12407 8472
rect 9673 8467 9739 8470
rect 12341 8467 12407 8470
rect 1761 8394 1827 8397
rect 18689 8394 18755 8397
rect 1761 8392 18755 8394
rect 1761 8336 1766 8392
rect 1822 8336 18694 8392
rect 18750 8336 18755 8392
rect 1761 8334 18755 8336
rect 1761 8331 1827 8334
rect 18689 8331 18755 8334
rect 0 8258 800 8288
rect 1393 8258 1459 8261
rect 0 8256 1459 8258
rect 0 8200 1398 8256
rect 1454 8200 1459 8256
rect 0 8198 1459 8200
rect 0 8168 800 8198
rect 1393 8195 1459 8198
rect 5576 8192 5896 8193
rect 5576 8128 5584 8192
rect 5648 8128 5664 8192
rect 5728 8128 5744 8192
rect 5808 8128 5824 8192
rect 5888 8128 5896 8192
rect 5576 8127 5896 8128
rect 14840 8192 15160 8193
rect 14840 8128 14848 8192
rect 14912 8128 14928 8192
rect 14992 8128 15008 8192
rect 15072 8128 15088 8192
rect 15152 8128 15160 8192
rect 14840 8127 15160 8128
rect 24104 8192 24424 8193
rect 24104 8128 24112 8192
rect 24176 8128 24192 8192
rect 24256 8128 24272 8192
rect 24336 8128 24352 8192
rect 24416 8128 24424 8192
rect 24104 8127 24424 8128
rect 10041 7986 10107 7989
rect 11094 7986 11100 7988
rect 10041 7984 11100 7986
rect 10041 7928 10046 7984
rect 10102 7928 11100 7984
rect 10041 7926 11100 7928
rect 10041 7923 10107 7926
rect 11094 7924 11100 7926
rect 11164 7924 11170 7988
rect 10208 7648 10528 7649
rect 10208 7584 10216 7648
rect 10280 7584 10296 7648
rect 10360 7584 10376 7648
rect 10440 7584 10456 7648
rect 10520 7584 10528 7648
rect 10208 7583 10528 7584
rect 19472 7648 19792 7649
rect 19472 7584 19480 7648
rect 19544 7584 19560 7648
rect 19624 7584 19640 7648
rect 19704 7584 19720 7648
rect 19784 7584 19792 7648
rect 19472 7583 19792 7584
rect 28349 7578 28415 7581
rect 29200 7578 30000 7608
rect 28349 7576 30000 7578
rect 28349 7520 28354 7576
rect 28410 7520 30000 7576
rect 28349 7518 30000 7520
rect 28349 7515 28415 7518
rect 29200 7488 30000 7518
rect 5576 7104 5896 7105
rect 5576 7040 5584 7104
rect 5648 7040 5664 7104
rect 5728 7040 5744 7104
rect 5808 7040 5824 7104
rect 5888 7040 5896 7104
rect 5576 7039 5896 7040
rect 14840 7104 15160 7105
rect 14840 7040 14848 7104
rect 14912 7040 14928 7104
rect 14992 7040 15008 7104
rect 15072 7040 15088 7104
rect 15152 7040 15160 7104
rect 14840 7039 15160 7040
rect 24104 7104 24424 7105
rect 24104 7040 24112 7104
rect 24176 7040 24192 7104
rect 24256 7040 24272 7104
rect 24336 7040 24352 7104
rect 24416 7040 24424 7104
rect 24104 7039 24424 7040
rect 0 6808 800 6928
rect 29200 6808 30000 6928
rect 10208 6560 10528 6561
rect 10208 6496 10216 6560
rect 10280 6496 10296 6560
rect 10360 6496 10376 6560
rect 10440 6496 10456 6560
rect 10520 6496 10528 6560
rect 10208 6495 10528 6496
rect 19472 6560 19792 6561
rect 19472 6496 19480 6560
rect 19544 6496 19560 6560
rect 19624 6496 19640 6560
rect 19704 6496 19720 6560
rect 19784 6496 19792 6560
rect 19472 6495 19792 6496
rect 5576 6016 5896 6017
rect 5576 5952 5584 6016
rect 5648 5952 5664 6016
rect 5728 5952 5744 6016
rect 5808 5952 5824 6016
rect 5888 5952 5896 6016
rect 5576 5951 5896 5952
rect 14840 6016 15160 6017
rect 14840 5952 14848 6016
rect 14912 5952 14928 6016
rect 14992 5952 15008 6016
rect 15072 5952 15088 6016
rect 15152 5952 15160 6016
rect 14840 5951 15160 5952
rect 24104 6016 24424 6017
rect 24104 5952 24112 6016
rect 24176 5952 24192 6016
rect 24256 5952 24272 6016
rect 24336 5952 24352 6016
rect 24416 5952 24424 6016
rect 24104 5951 24424 5952
rect 8477 5946 8543 5949
rect 14222 5946 14228 5948
rect 8477 5944 14228 5946
rect 8477 5888 8482 5944
rect 8538 5888 14228 5944
rect 8477 5886 14228 5888
rect 8477 5883 8543 5886
rect 14222 5884 14228 5886
rect 14292 5884 14298 5948
rect 10593 5674 10659 5677
rect 16573 5674 16639 5677
rect 10593 5672 16639 5674
rect 10593 5616 10598 5672
rect 10654 5616 16578 5672
rect 16634 5616 16639 5672
rect 10593 5614 16639 5616
rect 10593 5611 10659 5614
rect 16573 5611 16639 5614
rect 0 5538 800 5568
rect 1485 5538 1551 5541
rect 0 5536 1551 5538
rect 0 5480 1490 5536
rect 1546 5480 1551 5536
rect 0 5478 1551 5480
rect 0 5448 800 5478
rect 1485 5475 1551 5478
rect 28349 5538 28415 5541
rect 29200 5538 30000 5568
rect 28349 5536 30000 5538
rect 28349 5480 28354 5536
rect 28410 5480 30000 5536
rect 28349 5478 30000 5480
rect 28349 5475 28415 5478
rect 10208 5472 10528 5473
rect 10208 5408 10216 5472
rect 10280 5408 10296 5472
rect 10360 5408 10376 5472
rect 10440 5408 10456 5472
rect 10520 5408 10528 5472
rect 10208 5407 10528 5408
rect 19472 5472 19792 5473
rect 19472 5408 19480 5472
rect 19544 5408 19560 5472
rect 19624 5408 19640 5472
rect 19704 5408 19720 5472
rect 19784 5408 19792 5472
rect 29200 5448 30000 5478
rect 19472 5407 19792 5408
rect 12249 5130 12315 5133
rect 12249 5128 12450 5130
rect 12249 5072 12254 5128
rect 12310 5072 12450 5128
rect 12249 5070 12450 5072
rect 12249 5067 12315 5070
rect 12390 4994 12450 5070
rect 12525 4994 12591 4997
rect 12390 4992 12591 4994
rect 12390 4936 12530 4992
rect 12586 4936 12591 4992
rect 12390 4934 12591 4936
rect 12525 4931 12591 4934
rect 5576 4928 5896 4929
rect 5576 4864 5584 4928
rect 5648 4864 5664 4928
rect 5728 4864 5744 4928
rect 5808 4864 5824 4928
rect 5888 4864 5896 4928
rect 5576 4863 5896 4864
rect 14840 4928 15160 4929
rect 14840 4864 14848 4928
rect 14912 4864 14928 4928
rect 14992 4864 15008 4928
rect 15072 4864 15088 4928
rect 15152 4864 15160 4928
rect 14840 4863 15160 4864
rect 24104 4928 24424 4929
rect 24104 4864 24112 4928
rect 24176 4864 24192 4928
rect 24256 4864 24272 4928
rect 24336 4864 24352 4928
rect 24416 4864 24424 4928
rect 24104 4863 24424 4864
rect 10208 4384 10528 4385
rect 10208 4320 10216 4384
rect 10280 4320 10296 4384
rect 10360 4320 10376 4384
rect 10440 4320 10456 4384
rect 10520 4320 10528 4384
rect 10208 4319 10528 4320
rect 19472 4384 19792 4385
rect 19472 4320 19480 4384
rect 19544 4320 19560 4384
rect 19624 4320 19640 4384
rect 19704 4320 19720 4384
rect 19784 4320 19792 4384
rect 19472 4319 19792 4320
rect 0 4088 800 4208
rect 28349 4178 28415 4181
rect 29200 4178 30000 4208
rect 28349 4176 30000 4178
rect 28349 4120 28354 4176
rect 28410 4120 30000 4176
rect 28349 4118 30000 4120
rect 28349 4115 28415 4118
rect 29200 4088 30000 4118
rect 5576 3840 5896 3841
rect 5576 3776 5584 3840
rect 5648 3776 5664 3840
rect 5728 3776 5744 3840
rect 5808 3776 5824 3840
rect 5888 3776 5896 3840
rect 5576 3775 5896 3776
rect 14840 3840 15160 3841
rect 14840 3776 14848 3840
rect 14912 3776 14928 3840
rect 14992 3776 15008 3840
rect 15072 3776 15088 3840
rect 15152 3776 15160 3840
rect 14840 3775 15160 3776
rect 24104 3840 24424 3841
rect 24104 3776 24112 3840
rect 24176 3776 24192 3840
rect 24256 3776 24272 3840
rect 24336 3776 24352 3840
rect 24416 3776 24424 3840
rect 24104 3775 24424 3776
rect 0 3408 800 3528
rect 8201 3498 8267 3501
rect 13854 3498 13860 3500
rect 8201 3496 13860 3498
rect 8201 3440 8206 3496
rect 8262 3440 13860 3496
rect 8201 3438 13860 3440
rect 8201 3435 8267 3438
rect 13854 3436 13860 3438
rect 13924 3436 13930 3500
rect 29200 3408 30000 3528
rect 10208 3296 10528 3297
rect 10208 3232 10216 3296
rect 10280 3232 10296 3296
rect 10360 3232 10376 3296
rect 10440 3232 10456 3296
rect 10520 3232 10528 3296
rect 10208 3231 10528 3232
rect 19472 3296 19792 3297
rect 19472 3232 19480 3296
rect 19544 3232 19560 3296
rect 19624 3232 19640 3296
rect 19704 3232 19720 3296
rect 19784 3232 19792 3296
rect 19472 3231 19792 3232
rect 5576 2752 5896 2753
rect 5576 2688 5584 2752
rect 5648 2688 5664 2752
rect 5728 2688 5744 2752
rect 5808 2688 5824 2752
rect 5888 2688 5896 2752
rect 5576 2687 5896 2688
rect 14840 2752 15160 2753
rect 14840 2688 14848 2752
rect 14912 2688 14928 2752
rect 14992 2688 15008 2752
rect 15072 2688 15088 2752
rect 15152 2688 15160 2752
rect 14840 2687 15160 2688
rect 24104 2752 24424 2753
rect 24104 2688 24112 2752
rect 24176 2688 24192 2752
rect 24256 2688 24272 2752
rect 24336 2688 24352 2752
rect 24416 2688 24424 2752
rect 24104 2687 24424 2688
rect 10208 2208 10528 2209
rect 0 2138 800 2168
rect 10208 2144 10216 2208
rect 10280 2144 10296 2208
rect 10360 2144 10376 2208
rect 10440 2144 10456 2208
rect 10520 2144 10528 2208
rect 10208 2143 10528 2144
rect 19472 2208 19792 2209
rect 19472 2144 19480 2208
rect 19544 2144 19560 2208
rect 19624 2144 19640 2208
rect 19704 2144 19720 2208
rect 19784 2144 19792 2208
rect 19472 2143 19792 2144
rect 2221 2138 2287 2141
rect 0 2136 2287 2138
rect 0 2080 2226 2136
rect 2282 2080 2287 2136
rect 0 2078 2287 2080
rect 0 2048 800 2078
rect 2221 2075 2287 2078
rect 29200 2048 30000 2168
rect 0 778 800 808
rect 1669 778 1735 781
rect 0 776 1735 778
rect 0 720 1674 776
rect 1730 720 1735 776
rect 0 718 1735 720
rect 0 688 800 718
rect 1669 715 1735 718
rect 28257 778 28323 781
rect 29200 778 30000 808
rect 28257 776 30000 778
rect 28257 720 28262 776
rect 28318 720 30000 776
rect 28257 718 30000 720
rect 28257 715 28323 718
rect 29200 688 30000 718
<< via3 >>
rect 5584 27772 5648 27776
rect 5584 27716 5588 27772
rect 5588 27716 5644 27772
rect 5644 27716 5648 27772
rect 5584 27712 5648 27716
rect 5664 27772 5728 27776
rect 5664 27716 5668 27772
rect 5668 27716 5724 27772
rect 5724 27716 5728 27772
rect 5664 27712 5728 27716
rect 5744 27772 5808 27776
rect 5744 27716 5748 27772
rect 5748 27716 5804 27772
rect 5804 27716 5808 27772
rect 5744 27712 5808 27716
rect 5824 27772 5888 27776
rect 5824 27716 5828 27772
rect 5828 27716 5884 27772
rect 5884 27716 5888 27772
rect 5824 27712 5888 27716
rect 14848 27772 14912 27776
rect 14848 27716 14852 27772
rect 14852 27716 14908 27772
rect 14908 27716 14912 27772
rect 14848 27712 14912 27716
rect 14928 27772 14992 27776
rect 14928 27716 14932 27772
rect 14932 27716 14988 27772
rect 14988 27716 14992 27772
rect 14928 27712 14992 27716
rect 15008 27772 15072 27776
rect 15008 27716 15012 27772
rect 15012 27716 15068 27772
rect 15068 27716 15072 27772
rect 15008 27712 15072 27716
rect 15088 27772 15152 27776
rect 15088 27716 15092 27772
rect 15092 27716 15148 27772
rect 15148 27716 15152 27772
rect 15088 27712 15152 27716
rect 24112 27772 24176 27776
rect 24112 27716 24116 27772
rect 24116 27716 24172 27772
rect 24172 27716 24176 27772
rect 24112 27712 24176 27716
rect 24192 27772 24256 27776
rect 24192 27716 24196 27772
rect 24196 27716 24252 27772
rect 24252 27716 24256 27772
rect 24192 27712 24256 27716
rect 24272 27772 24336 27776
rect 24272 27716 24276 27772
rect 24276 27716 24332 27772
rect 24332 27716 24336 27772
rect 24272 27712 24336 27716
rect 24352 27772 24416 27776
rect 24352 27716 24356 27772
rect 24356 27716 24412 27772
rect 24412 27716 24416 27772
rect 24352 27712 24416 27716
rect 10216 27228 10280 27232
rect 10216 27172 10220 27228
rect 10220 27172 10276 27228
rect 10276 27172 10280 27228
rect 10216 27168 10280 27172
rect 10296 27228 10360 27232
rect 10296 27172 10300 27228
rect 10300 27172 10356 27228
rect 10356 27172 10360 27228
rect 10296 27168 10360 27172
rect 10376 27228 10440 27232
rect 10376 27172 10380 27228
rect 10380 27172 10436 27228
rect 10436 27172 10440 27228
rect 10376 27168 10440 27172
rect 10456 27228 10520 27232
rect 10456 27172 10460 27228
rect 10460 27172 10516 27228
rect 10516 27172 10520 27228
rect 10456 27168 10520 27172
rect 19480 27228 19544 27232
rect 19480 27172 19484 27228
rect 19484 27172 19540 27228
rect 19540 27172 19544 27228
rect 19480 27168 19544 27172
rect 19560 27228 19624 27232
rect 19560 27172 19564 27228
rect 19564 27172 19620 27228
rect 19620 27172 19624 27228
rect 19560 27168 19624 27172
rect 19640 27228 19704 27232
rect 19640 27172 19644 27228
rect 19644 27172 19700 27228
rect 19700 27172 19704 27228
rect 19640 27168 19704 27172
rect 19720 27228 19784 27232
rect 19720 27172 19724 27228
rect 19724 27172 19780 27228
rect 19780 27172 19784 27228
rect 19720 27168 19784 27172
rect 5584 26684 5648 26688
rect 5584 26628 5588 26684
rect 5588 26628 5644 26684
rect 5644 26628 5648 26684
rect 5584 26624 5648 26628
rect 5664 26684 5728 26688
rect 5664 26628 5668 26684
rect 5668 26628 5724 26684
rect 5724 26628 5728 26684
rect 5664 26624 5728 26628
rect 5744 26684 5808 26688
rect 5744 26628 5748 26684
rect 5748 26628 5804 26684
rect 5804 26628 5808 26684
rect 5744 26624 5808 26628
rect 5824 26684 5888 26688
rect 5824 26628 5828 26684
rect 5828 26628 5884 26684
rect 5884 26628 5888 26684
rect 5824 26624 5888 26628
rect 14848 26684 14912 26688
rect 14848 26628 14852 26684
rect 14852 26628 14908 26684
rect 14908 26628 14912 26684
rect 14848 26624 14912 26628
rect 14928 26684 14992 26688
rect 14928 26628 14932 26684
rect 14932 26628 14988 26684
rect 14988 26628 14992 26684
rect 14928 26624 14992 26628
rect 15008 26684 15072 26688
rect 15008 26628 15012 26684
rect 15012 26628 15068 26684
rect 15068 26628 15072 26684
rect 15008 26624 15072 26628
rect 15088 26684 15152 26688
rect 15088 26628 15092 26684
rect 15092 26628 15148 26684
rect 15148 26628 15152 26684
rect 15088 26624 15152 26628
rect 24112 26684 24176 26688
rect 24112 26628 24116 26684
rect 24116 26628 24172 26684
rect 24172 26628 24176 26684
rect 24112 26624 24176 26628
rect 24192 26684 24256 26688
rect 24192 26628 24196 26684
rect 24196 26628 24252 26684
rect 24252 26628 24256 26684
rect 24192 26624 24256 26628
rect 24272 26684 24336 26688
rect 24272 26628 24276 26684
rect 24276 26628 24332 26684
rect 24332 26628 24336 26684
rect 24272 26624 24336 26628
rect 24352 26684 24416 26688
rect 24352 26628 24356 26684
rect 24356 26628 24412 26684
rect 24412 26628 24416 26684
rect 24352 26624 24416 26628
rect 10216 26140 10280 26144
rect 10216 26084 10220 26140
rect 10220 26084 10276 26140
rect 10276 26084 10280 26140
rect 10216 26080 10280 26084
rect 10296 26140 10360 26144
rect 10296 26084 10300 26140
rect 10300 26084 10356 26140
rect 10356 26084 10360 26140
rect 10296 26080 10360 26084
rect 10376 26140 10440 26144
rect 10376 26084 10380 26140
rect 10380 26084 10436 26140
rect 10436 26084 10440 26140
rect 10376 26080 10440 26084
rect 10456 26140 10520 26144
rect 10456 26084 10460 26140
rect 10460 26084 10516 26140
rect 10516 26084 10520 26140
rect 10456 26080 10520 26084
rect 19480 26140 19544 26144
rect 19480 26084 19484 26140
rect 19484 26084 19540 26140
rect 19540 26084 19544 26140
rect 19480 26080 19544 26084
rect 19560 26140 19624 26144
rect 19560 26084 19564 26140
rect 19564 26084 19620 26140
rect 19620 26084 19624 26140
rect 19560 26080 19624 26084
rect 19640 26140 19704 26144
rect 19640 26084 19644 26140
rect 19644 26084 19700 26140
rect 19700 26084 19704 26140
rect 19640 26080 19704 26084
rect 19720 26140 19784 26144
rect 19720 26084 19724 26140
rect 19724 26084 19780 26140
rect 19780 26084 19784 26140
rect 19720 26080 19784 26084
rect 5584 25596 5648 25600
rect 5584 25540 5588 25596
rect 5588 25540 5644 25596
rect 5644 25540 5648 25596
rect 5584 25536 5648 25540
rect 5664 25596 5728 25600
rect 5664 25540 5668 25596
rect 5668 25540 5724 25596
rect 5724 25540 5728 25596
rect 5664 25536 5728 25540
rect 5744 25596 5808 25600
rect 5744 25540 5748 25596
rect 5748 25540 5804 25596
rect 5804 25540 5808 25596
rect 5744 25536 5808 25540
rect 5824 25596 5888 25600
rect 5824 25540 5828 25596
rect 5828 25540 5884 25596
rect 5884 25540 5888 25596
rect 5824 25536 5888 25540
rect 14848 25596 14912 25600
rect 14848 25540 14852 25596
rect 14852 25540 14908 25596
rect 14908 25540 14912 25596
rect 14848 25536 14912 25540
rect 14928 25596 14992 25600
rect 14928 25540 14932 25596
rect 14932 25540 14988 25596
rect 14988 25540 14992 25596
rect 14928 25536 14992 25540
rect 15008 25596 15072 25600
rect 15008 25540 15012 25596
rect 15012 25540 15068 25596
rect 15068 25540 15072 25596
rect 15008 25536 15072 25540
rect 15088 25596 15152 25600
rect 15088 25540 15092 25596
rect 15092 25540 15148 25596
rect 15148 25540 15152 25596
rect 15088 25536 15152 25540
rect 24112 25596 24176 25600
rect 24112 25540 24116 25596
rect 24116 25540 24172 25596
rect 24172 25540 24176 25596
rect 24112 25536 24176 25540
rect 24192 25596 24256 25600
rect 24192 25540 24196 25596
rect 24196 25540 24252 25596
rect 24252 25540 24256 25596
rect 24192 25536 24256 25540
rect 24272 25596 24336 25600
rect 24272 25540 24276 25596
rect 24276 25540 24332 25596
rect 24332 25540 24336 25596
rect 24272 25536 24336 25540
rect 24352 25596 24416 25600
rect 24352 25540 24356 25596
rect 24356 25540 24412 25596
rect 24412 25540 24416 25596
rect 24352 25536 24416 25540
rect 10216 25052 10280 25056
rect 10216 24996 10220 25052
rect 10220 24996 10276 25052
rect 10276 24996 10280 25052
rect 10216 24992 10280 24996
rect 10296 25052 10360 25056
rect 10296 24996 10300 25052
rect 10300 24996 10356 25052
rect 10356 24996 10360 25052
rect 10296 24992 10360 24996
rect 10376 25052 10440 25056
rect 10376 24996 10380 25052
rect 10380 24996 10436 25052
rect 10436 24996 10440 25052
rect 10376 24992 10440 24996
rect 10456 25052 10520 25056
rect 10456 24996 10460 25052
rect 10460 24996 10516 25052
rect 10516 24996 10520 25052
rect 10456 24992 10520 24996
rect 19480 25052 19544 25056
rect 19480 24996 19484 25052
rect 19484 24996 19540 25052
rect 19540 24996 19544 25052
rect 19480 24992 19544 24996
rect 19560 25052 19624 25056
rect 19560 24996 19564 25052
rect 19564 24996 19620 25052
rect 19620 24996 19624 25052
rect 19560 24992 19624 24996
rect 19640 25052 19704 25056
rect 19640 24996 19644 25052
rect 19644 24996 19700 25052
rect 19700 24996 19704 25052
rect 19640 24992 19704 24996
rect 19720 25052 19784 25056
rect 19720 24996 19724 25052
rect 19724 24996 19780 25052
rect 19780 24996 19784 25052
rect 19720 24992 19784 24996
rect 5584 24508 5648 24512
rect 5584 24452 5588 24508
rect 5588 24452 5644 24508
rect 5644 24452 5648 24508
rect 5584 24448 5648 24452
rect 5664 24508 5728 24512
rect 5664 24452 5668 24508
rect 5668 24452 5724 24508
rect 5724 24452 5728 24508
rect 5664 24448 5728 24452
rect 5744 24508 5808 24512
rect 5744 24452 5748 24508
rect 5748 24452 5804 24508
rect 5804 24452 5808 24508
rect 5744 24448 5808 24452
rect 5824 24508 5888 24512
rect 5824 24452 5828 24508
rect 5828 24452 5884 24508
rect 5884 24452 5888 24508
rect 5824 24448 5888 24452
rect 14848 24508 14912 24512
rect 14848 24452 14852 24508
rect 14852 24452 14908 24508
rect 14908 24452 14912 24508
rect 14848 24448 14912 24452
rect 14928 24508 14992 24512
rect 14928 24452 14932 24508
rect 14932 24452 14988 24508
rect 14988 24452 14992 24508
rect 14928 24448 14992 24452
rect 15008 24508 15072 24512
rect 15008 24452 15012 24508
rect 15012 24452 15068 24508
rect 15068 24452 15072 24508
rect 15008 24448 15072 24452
rect 15088 24508 15152 24512
rect 15088 24452 15092 24508
rect 15092 24452 15148 24508
rect 15148 24452 15152 24508
rect 15088 24448 15152 24452
rect 24112 24508 24176 24512
rect 24112 24452 24116 24508
rect 24116 24452 24172 24508
rect 24172 24452 24176 24508
rect 24112 24448 24176 24452
rect 24192 24508 24256 24512
rect 24192 24452 24196 24508
rect 24196 24452 24252 24508
rect 24252 24452 24256 24508
rect 24192 24448 24256 24452
rect 24272 24508 24336 24512
rect 24272 24452 24276 24508
rect 24276 24452 24332 24508
rect 24332 24452 24336 24508
rect 24272 24448 24336 24452
rect 24352 24508 24416 24512
rect 24352 24452 24356 24508
rect 24356 24452 24412 24508
rect 24412 24452 24416 24508
rect 24352 24448 24416 24452
rect 10216 23964 10280 23968
rect 10216 23908 10220 23964
rect 10220 23908 10276 23964
rect 10276 23908 10280 23964
rect 10216 23904 10280 23908
rect 10296 23964 10360 23968
rect 10296 23908 10300 23964
rect 10300 23908 10356 23964
rect 10356 23908 10360 23964
rect 10296 23904 10360 23908
rect 10376 23964 10440 23968
rect 10376 23908 10380 23964
rect 10380 23908 10436 23964
rect 10436 23908 10440 23964
rect 10376 23904 10440 23908
rect 10456 23964 10520 23968
rect 10456 23908 10460 23964
rect 10460 23908 10516 23964
rect 10516 23908 10520 23964
rect 10456 23904 10520 23908
rect 19480 23964 19544 23968
rect 19480 23908 19484 23964
rect 19484 23908 19540 23964
rect 19540 23908 19544 23964
rect 19480 23904 19544 23908
rect 19560 23964 19624 23968
rect 19560 23908 19564 23964
rect 19564 23908 19620 23964
rect 19620 23908 19624 23964
rect 19560 23904 19624 23908
rect 19640 23964 19704 23968
rect 19640 23908 19644 23964
rect 19644 23908 19700 23964
rect 19700 23908 19704 23964
rect 19640 23904 19704 23908
rect 19720 23964 19784 23968
rect 19720 23908 19724 23964
rect 19724 23908 19780 23964
rect 19780 23908 19784 23964
rect 19720 23904 19784 23908
rect 5584 23420 5648 23424
rect 5584 23364 5588 23420
rect 5588 23364 5644 23420
rect 5644 23364 5648 23420
rect 5584 23360 5648 23364
rect 5664 23420 5728 23424
rect 5664 23364 5668 23420
rect 5668 23364 5724 23420
rect 5724 23364 5728 23420
rect 5664 23360 5728 23364
rect 5744 23420 5808 23424
rect 5744 23364 5748 23420
rect 5748 23364 5804 23420
rect 5804 23364 5808 23420
rect 5744 23360 5808 23364
rect 5824 23420 5888 23424
rect 5824 23364 5828 23420
rect 5828 23364 5884 23420
rect 5884 23364 5888 23420
rect 5824 23360 5888 23364
rect 14848 23420 14912 23424
rect 14848 23364 14852 23420
rect 14852 23364 14908 23420
rect 14908 23364 14912 23420
rect 14848 23360 14912 23364
rect 14928 23420 14992 23424
rect 14928 23364 14932 23420
rect 14932 23364 14988 23420
rect 14988 23364 14992 23420
rect 14928 23360 14992 23364
rect 15008 23420 15072 23424
rect 15008 23364 15012 23420
rect 15012 23364 15068 23420
rect 15068 23364 15072 23420
rect 15008 23360 15072 23364
rect 15088 23420 15152 23424
rect 15088 23364 15092 23420
rect 15092 23364 15148 23420
rect 15148 23364 15152 23420
rect 15088 23360 15152 23364
rect 24112 23420 24176 23424
rect 24112 23364 24116 23420
rect 24116 23364 24172 23420
rect 24172 23364 24176 23420
rect 24112 23360 24176 23364
rect 24192 23420 24256 23424
rect 24192 23364 24196 23420
rect 24196 23364 24252 23420
rect 24252 23364 24256 23420
rect 24192 23360 24256 23364
rect 24272 23420 24336 23424
rect 24272 23364 24276 23420
rect 24276 23364 24332 23420
rect 24332 23364 24336 23420
rect 24272 23360 24336 23364
rect 24352 23420 24416 23424
rect 24352 23364 24356 23420
rect 24356 23364 24412 23420
rect 24412 23364 24416 23420
rect 24352 23360 24416 23364
rect 10216 22876 10280 22880
rect 10216 22820 10220 22876
rect 10220 22820 10276 22876
rect 10276 22820 10280 22876
rect 10216 22816 10280 22820
rect 10296 22876 10360 22880
rect 10296 22820 10300 22876
rect 10300 22820 10356 22876
rect 10356 22820 10360 22876
rect 10296 22816 10360 22820
rect 10376 22876 10440 22880
rect 10376 22820 10380 22876
rect 10380 22820 10436 22876
rect 10436 22820 10440 22876
rect 10376 22816 10440 22820
rect 10456 22876 10520 22880
rect 10456 22820 10460 22876
rect 10460 22820 10516 22876
rect 10516 22820 10520 22876
rect 10456 22816 10520 22820
rect 19480 22876 19544 22880
rect 19480 22820 19484 22876
rect 19484 22820 19540 22876
rect 19540 22820 19544 22876
rect 19480 22816 19544 22820
rect 19560 22876 19624 22880
rect 19560 22820 19564 22876
rect 19564 22820 19620 22876
rect 19620 22820 19624 22876
rect 19560 22816 19624 22820
rect 19640 22876 19704 22880
rect 19640 22820 19644 22876
rect 19644 22820 19700 22876
rect 19700 22820 19704 22876
rect 19640 22816 19704 22820
rect 19720 22876 19784 22880
rect 19720 22820 19724 22876
rect 19724 22820 19780 22876
rect 19780 22820 19784 22876
rect 19720 22816 19784 22820
rect 5584 22332 5648 22336
rect 5584 22276 5588 22332
rect 5588 22276 5644 22332
rect 5644 22276 5648 22332
rect 5584 22272 5648 22276
rect 5664 22332 5728 22336
rect 5664 22276 5668 22332
rect 5668 22276 5724 22332
rect 5724 22276 5728 22332
rect 5664 22272 5728 22276
rect 5744 22332 5808 22336
rect 5744 22276 5748 22332
rect 5748 22276 5804 22332
rect 5804 22276 5808 22332
rect 5744 22272 5808 22276
rect 5824 22332 5888 22336
rect 5824 22276 5828 22332
rect 5828 22276 5884 22332
rect 5884 22276 5888 22332
rect 5824 22272 5888 22276
rect 14848 22332 14912 22336
rect 14848 22276 14852 22332
rect 14852 22276 14908 22332
rect 14908 22276 14912 22332
rect 14848 22272 14912 22276
rect 14928 22332 14992 22336
rect 14928 22276 14932 22332
rect 14932 22276 14988 22332
rect 14988 22276 14992 22332
rect 14928 22272 14992 22276
rect 15008 22332 15072 22336
rect 15008 22276 15012 22332
rect 15012 22276 15068 22332
rect 15068 22276 15072 22332
rect 15008 22272 15072 22276
rect 15088 22332 15152 22336
rect 15088 22276 15092 22332
rect 15092 22276 15148 22332
rect 15148 22276 15152 22332
rect 15088 22272 15152 22276
rect 24112 22332 24176 22336
rect 24112 22276 24116 22332
rect 24116 22276 24172 22332
rect 24172 22276 24176 22332
rect 24112 22272 24176 22276
rect 24192 22332 24256 22336
rect 24192 22276 24196 22332
rect 24196 22276 24252 22332
rect 24252 22276 24256 22332
rect 24192 22272 24256 22276
rect 24272 22332 24336 22336
rect 24272 22276 24276 22332
rect 24276 22276 24332 22332
rect 24332 22276 24336 22332
rect 24272 22272 24336 22276
rect 24352 22332 24416 22336
rect 24352 22276 24356 22332
rect 24356 22276 24412 22332
rect 24412 22276 24416 22332
rect 24352 22272 24416 22276
rect 10216 21788 10280 21792
rect 10216 21732 10220 21788
rect 10220 21732 10276 21788
rect 10276 21732 10280 21788
rect 10216 21728 10280 21732
rect 10296 21788 10360 21792
rect 10296 21732 10300 21788
rect 10300 21732 10356 21788
rect 10356 21732 10360 21788
rect 10296 21728 10360 21732
rect 10376 21788 10440 21792
rect 10376 21732 10380 21788
rect 10380 21732 10436 21788
rect 10436 21732 10440 21788
rect 10376 21728 10440 21732
rect 10456 21788 10520 21792
rect 10456 21732 10460 21788
rect 10460 21732 10516 21788
rect 10516 21732 10520 21788
rect 10456 21728 10520 21732
rect 19480 21788 19544 21792
rect 19480 21732 19484 21788
rect 19484 21732 19540 21788
rect 19540 21732 19544 21788
rect 19480 21728 19544 21732
rect 19560 21788 19624 21792
rect 19560 21732 19564 21788
rect 19564 21732 19620 21788
rect 19620 21732 19624 21788
rect 19560 21728 19624 21732
rect 19640 21788 19704 21792
rect 19640 21732 19644 21788
rect 19644 21732 19700 21788
rect 19700 21732 19704 21788
rect 19640 21728 19704 21732
rect 19720 21788 19784 21792
rect 19720 21732 19724 21788
rect 19724 21732 19780 21788
rect 19780 21732 19784 21788
rect 19720 21728 19784 21732
rect 17540 21252 17604 21316
rect 5584 21244 5648 21248
rect 5584 21188 5588 21244
rect 5588 21188 5644 21244
rect 5644 21188 5648 21244
rect 5584 21184 5648 21188
rect 5664 21244 5728 21248
rect 5664 21188 5668 21244
rect 5668 21188 5724 21244
rect 5724 21188 5728 21244
rect 5664 21184 5728 21188
rect 5744 21244 5808 21248
rect 5744 21188 5748 21244
rect 5748 21188 5804 21244
rect 5804 21188 5808 21244
rect 5744 21184 5808 21188
rect 5824 21244 5888 21248
rect 5824 21188 5828 21244
rect 5828 21188 5884 21244
rect 5884 21188 5888 21244
rect 5824 21184 5888 21188
rect 14848 21244 14912 21248
rect 14848 21188 14852 21244
rect 14852 21188 14908 21244
rect 14908 21188 14912 21244
rect 14848 21184 14912 21188
rect 14928 21244 14992 21248
rect 14928 21188 14932 21244
rect 14932 21188 14988 21244
rect 14988 21188 14992 21244
rect 14928 21184 14992 21188
rect 15008 21244 15072 21248
rect 15008 21188 15012 21244
rect 15012 21188 15068 21244
rect 15068 21188 15072 21244
rect 15008 21184 15072 21188
rect 15088 21244 15152 21248
rect 15088 21188 15092 21244
rect 15092 21188 15148 21244
rect 15148 21188 15152 21244
rect 15088 21184 15152 21188
rect 24112 21244 24176 21248
rect 24112 21188 24116 21244
rect 24116 21188 24172 21244
rect 24172 21188 24176 21244
rect 24112 21184 24176 21188
rect 24192 21244 24256 21248
rect 24192 21188 24196 21244
rect 24196 21188 24252 21244
rect 24252 21188 24256 21244
rect 24192 21184 24256 21188
rect 24272 21244 24336 21248
rect 24272 21188 24276 21244
rect 24276 21188 24332 21244
rect 24332 21188 24336 21244
rect 24272 21184 24336 21188
rect 24352 21244 24416 21248
rect 24352 21188 24356 21244
rect 24356 21188 24412 21244
rect 24412 21188 24416 21244
rect 24352 21184 24416 21188
rect 10216 20700 10280 20704
rect 10216 20644 10220 20700
rect 10220 20644 10276 20700
rect 10276 20644 10280 20700
rect 10216 20640 10280 20644
rect 10296 20700 10360 20704
rect 10296 20644 10300 20700
rect 10300 20644 10356 20700
rect 10356 20644 10360 20700
rect 10296 20640 10360 20644
rect 10376 20700 10440 20704
rect 10376 20644 10380 20700
rect 10380 20644 10436 20700
rect 10436 20644 10440 20700
rect 10376 20640 10440 20644
rect 10456 20700 10520 20704
rect 10456 20644 10460 20700
rect 10460 20644 10516 20700
rect 10516 20644 10520 20700
rect 10456 20640 10520 20644
rect 19480 20700 19544 20704
rect 19480 20644 19484 20700
rect 19484 20644 19540 20700
rect 19540 20644 19544 20700
rect 19480 20640 19544 20644
rect 19560 20700 19624 20704
rect 19560 20644 19564 20700
rect 19564 20644 19620 20700
rect 19620 20644 19624 20700
rect 19560 20640 19624 20644
rect 19640 20700 19704 20704
rect 19640 20644 19644 20700
rect 19644 20644 19700 20700
rect 19700 20644 19704 20700
rect 19640 20640 19704 20644
rect 19720 20700 19784 20704
rect 19720 20644 19724 20700
rect 19724 20644 19780 20700
rect 19780 20644 19784 20700
rect 19720 20640 19784 20644
rect 5584 20156 5648 20160
rect 5584 20100 5588 20156
rect 5588 20100 5644 20156
rect 5644 20100 5648 20156
rect 5584 20096 5648 20100
rect 5664 20156 5728 20160
rect 5664 20100 5668 20156
rect 5668 20100 5724 20156
rect 5724 20100 5728 20156
rect 5664 20096 5728 20100
rect 5744 20156 5808 20160
rect 5744 20100 5748 20156
rect 5748 20100 5804 20156
rect 5804 20100 5808 20156
rect 5744 20096 5808 20100
rect 5824 20156 5888 20160
rect 5824 20100 5828 20156
rect 5828 20100 5884 20156
rect 5884 20100 5888 20156
rect 5824 20096 5888 20100
rect 14848 20156 14912 20160
rect 14848 20100 14852 20156
rect 14852 20100 14908 20156
rect 14908 20100 14912 20156
rect 14848 20096 14912 20100
rect 14928 20156 14992 20160
rect 14928 20100 14932 20156
rect 14932 20100 14988 20156
rect 14988 20100 14992 20156
rect 14928 20096 14992 20100
rect 15008 20156 15072 20160
rect 15008 20100 15012 20156
rect 15012 20100 15068 20156
rect 15068 20100 15072 20156
rect 15008 20096 15072 20100
rect 15088 20156 15152 20160
rect 15088 20100 15092 20156
rect 15092 20100 15148 20156
rect 15148 20100 15152 20156
rect 15088 20096 15152 20100
rect 24112 20156 24176 20160
rect 24112 20100 24116 20156
rect 24116 20100 24172 20156
rect 24172 20100 24176 20156
rect 24112 20096 24176 20100
rect 24192 20156 24256 20160
rect 24192 20100 24196 20156
rect 24196 20100 24252 20156
rect 24252 20100 24256 20156
rect 24192 20096 24256 20100
rect 24272 20156 24336 20160
rect 24272 20100 24276 20156
rect 24276 20100 24332 20156
rect 24332 20100 24336 20156
rect 24272 20096 24336 20100
rect 24352 20156 24416 20160
rect 24352 20100 24356 20156
rect 24356 20100 24412 20156
rect 24412 20100 24416 20156
rect 24352 20096 24416 20100
rect 21036 19680 21100 19684
rect 21036 19624 21086 19680
rect 21086 19624 21100 19680
rect 21036 19620 21100 19624
rect 10216 19612 10280 19616
rect 10216 19556 10220 19612
rect 10220 19556 10276 19612
rect 10276 19556 10280 19612
rect 10216 19552 10280 19556
rect 10296 19612 10360 19616
rect 10296 19556 10300 19612
rect 10300 19556 10356 19612
rect 10356 19556 10360 19612
rect 10296 19552 10360 19556
rect 10376 19612 10440 19616
rect 10376 19556 10380 19612
rect 10380 19556 10436 19612
rect 10436 19556 10440 19612
rect 10376 19552 10440 19556
rect 10456 19612 10520 19616
rect 10456 19556 10460 19612
rect 10460 19556 10516 19612
rect 10516 19556 10520 19612
rect 10456 19552 10520 19556
rect 19480 19612 19544 19616
rect 19480 19556 19484 19612
rect 19484 19556 19540 19612
rect 19540 19556 19544 19612
rect 19480 19552 19544 19556
rect 19560 19612 19624 19616
rect 19560 19556 19564 19612
rect 19564 19556 19620 19612
rect 19620 19556 19624 19612
rect 19560 19552 19624 19556
rect 19640 19612 19704 19616
rect 19640 19556 19644 19612
rect 19644 19556 19700 19612
rect 19700 19556 19704 19612
rect 19640 19552 19704 19556
rect 19720 19612 19784 19616
rect 19720 19556 19724 19612
rect 19724 19556 19780 19612
rect 19780 19556 19784 19612
rect 19720 19552 19784 19556
rect 5584 19068 5648 19072
rect 5584 19012 5588 19068
rect 5588 19012 5644 19068
rect 5644 19012 5648 19068
rect 5584 19008 5648 19012
rect 5664 19068 5728 19072
rect 5664 19012 5668 19068
rect 5668 19012 5724 19068
rect 5724 19012 5728 19068
rect 5664 19008 5728 19012
rect 5744 19068 5808 19072
rect 5744 19012 5748 19068
rect 5748 19012 5804 19068
rect 5804 19012 5808 19068
rect 5744 19008 5808 19012
rect 5824 19068 5888 19072
rect 5824 19012 5828 19068
rect 5828 19012 5884 19068
rect 5884 19012 5888 19068
rect 5824 19008 5888 19012
rect 14848 19068 14912 19072
rect 14848 19012 14852 19068
rect 14852 19012 14908 19068
rect 14908 19012 14912 19068
rect 14848 19008 14912 19012
rect 14928 19068 14992 19072
rect 14928 19012 14932 19068
rect 14932 19012 14988 19068
rect 14988 19012 14992 19068
rect 14928 19008 14992 19012
rect 15008 19068 15072 19072
rect 15008 19012 15012 19068
rect 15012 19012 15068 19068
rect 15068 19012 15072 19068
rect 15008 19008 15072 19012
rect 15088 19068 15152 19072
rect 15088 19012 15092 19068
rect 15092 19012 15148 19068
rect 15148 19012 15152 19068
rect 15088 19008 15152 19012
rect 24112 19068 24176 19072
rect 24112 19012 24116 19068
rect 24116 19012 24172 19068
rect 24172 19012 24176 19068
rect 24112 19008 24176 19012
rect 24192 19068 24256 19072
rect 24192 19012 24196 19068
rect 24196 19012 24252 19068
rect 24252 19012 24256 19068
rect 24192 19008 24256 19012
rect 24272 19068 24336 19072
rect 24272 19012 24276 19068
rect 24276 19012 24332 19068
rect 24332 19012 24336 19068
rect 24272 19008 24336 19012
rect 24352 19068 24416 19072
rect 24352 19012 24356 19068
rect 24356 19012 24412 19068
rect 24412 19012 24416 19068
rect 24352 19008 24416 19012
rect 10216 18524 10280 18528
rect 10216 18468 10220 18524
rect 10220 18468 10276 18524
rect 10276 18468 10280 18524
rect 10216 18464 10280 18468
rect 10296 18524 10360 18528
rect 10296 18468 10300 18524
rect 10300 18468 10356 18524
rect 10356 18468 10360 18524
rect 10296 18464 10360 18468
rect 10376 18524 10440 18528
rect 10376 18468 10380 18524
rect 10380 18468 10436 18524
rect 10436 18468 10440 18524
rect 10376 18464 10440 18468
rect 10456 18524 10520 18528
rect 10456 18468 10460 18524
rect 10460 18468 10516 18524
rect 10516 18468 10520 18524
rect 10456 18464 10520 18468
rect 19480 18524 19544 18528
rect 19480 18468 19484 18524
rect 19484 18468 19540 18524
rect 19540 18468 19544 18524
rect 19480 18464 19544 18468
rect 19560 18524 19624 18528
rect 19560 18468 19564 18524
rect 19564 18468 19620 18524
rect 19620 18468 19624 18524
rect 19560 18464 19624 18468
rect 19640 18524 19704 18528
rect 19640 18468 19644 18524
rect 19644 18468 19700 18524
rect 19700 18468 19704 18524
rect 19640 18464 19704 18468
rect 19720 18524 19784 18528
rect 19720 18468 19724 18524
rect 19724 18468 19780 18524
rect 19780 18468 19784 18524
rect 19720 18464 19784 18468
rect 5584 17980 5648 17984
rect 5584 17924 5588 17980
rect 5588 17924 5644 17980
rect 5644 17924 5648 17980
rect 5584 17920 5648 17924
rect 5664 17980 5728 17984
rect 5664 17924 5668 17980
rect 5668 17924 5724 17980
rect 5724 17924 5728 17980
rect 5664 17920 5728 17924
rect 5744 17980 5808 17984
rect 5744 17924 5748 17980
rect 5748 17924 5804 17980
rect 5804 17924 5808 17980
rect 5744 17920 5808 17924
rect 5824 17980 5888 17984
rect 5824 17924 5828 17980
rect 5828 17924 5884 17980
rect 5884 17924 5888 17980
rect 5824 17920 5888 17924
rect 14848 17980 14912 17984
rect 14848 17924 14852 17980
rect 14852 17924 14908 17980
rect 14908 17924 14912 17980
rect 14848 17920 14912 17924
rect 14928 17980 14992 17984
rect 14928 17924 14932 17980
rect 14932 17924 14988 17980
rect 14988 17924 14992 17980
rect 14928 17920 14992 17924
rect 15008 17980 15072 17984
rect 15008 17924 15012 17980
rect 15012 17924 15068 17980
rect 15068 17924 15072 17980
rect 15008 17920 15072 17924
rect 15088 17980 15152 17984
rect 15088 17924 15092 17980
rect 15092 17924 15148 17980
rect 15148 17924 15152 17980
rect 15088 17920 15152 17924
rect 24112 17980 24176 17984
rect 24112 17924 24116 17980
rect 24116 17924 24172 17980
rect 24172 17924 24176 17980
rect 24112 17920 24176 17924
rect 24192 17980 24256 17984
rect 24192 17924 24196 17980
rect 24196 17924 24252 17980
rect 24252 17924 24256 17980
rect 24192 17920 24256 17924
rect 24272 17980 24336 17984
rect 24272 17924 24276 17980
rect 24276 17924 24332 17980
rect 24332 17924 24336 17980
rect 24272 17920 24336 17924
rect 24352 17980 24416 17984
rect 24352 17924 24356 17980
rect 24356 17924 24412 17980
rect 24412 17924 24416 17980
rect 24352 17920 24416 17924
rect 10216 17436 10280 17440
rect 10216 17380 10220 17436
rect 10220 17380 10276 17436
rect 10276 17380 10280 17436
rect 10216 17376 10280 17380
rect 10296 17436 10360 17440
rect 10296 17380 10300 17436
rect 10300 17380 10356 17436
rect 10356 17380 10360 17436
rect 10296 17376 10360 17380
rect 10376 17436 10440 17440
rect 10376 17380 10380 17436
rect 10380 17380 10436 17436
rect 10436 17380 10440 17436
rect 10376 17376 10440 17380
rect 10456 17436 10520 17440
rect 10456 17380 10460 17436
rect 10460 17380 10516 17436
rect 10516 17380 10520 17436
rect 10456 17376 10520 17380
rect 19480 17436 19544 17440
rect 19480 17380 19484 17436
rect 19484 17380 19540 17436
rect 19540 17380 19544 17436
rect 19480 17376 19544 17380
rect 19560 17436 19624 17440
rect 19560 17380 19564 17436
rect 19564 17380 19620 17436
rect 19620 17380 19624 17436
rect 19560 17376 19624 17380
rect 19640 17436 19704 17440
rect 19640 17380 19644 17436
rect 19644 17380 19700 17436
rect 19700 17380 19704 17436
rect 19640 17376 19704 17380
rect 19720 17436 19784 17440
rect 19720 17380 19724 17436
rect 19724 17380 19780 17436
rect 19780 17380 19784 17436
rect 19720 17376 19784 17380
rect 5584 16892 5648 16896
rect 5584 16836 5588 16892
rect 5588 16836 5644 16892
rect 5644 16836 5648 16892
rect 5584 16832 5648 16836
rect 5664 16892 5728 16896
rect 5664 16836 5668 16892
rect 5668 16836 5724 16892
rect 5724 16836 5728 16892
rect 5664 16832 5728 16836
rect 5744 16892 5808 16896
rect 5744 16836 5748 16892
rect 5748 16836 5804 16892
rect 5804 16836 5808 16892
rect 5744 16832 5808 16836
rect 5824 16892 5888 16896
rect 5824 16836 5828 16892
rect 5828 16836 5884 16892
rect 5884 16836 5888 16892
rect 5824 16832 5888 16836
rect 14848 16892 14912 16896
rect 14848 16836 14852 16892
rect 14852 16836 14908 16892
rect 14908 16836 14912 16892
rect 14848 16832 14912 16836
rect 14928 16892 14992 16896
rect 14928 16836 14932 16892
rect 14932 16836 14988 16892
rect 14988 16836 14992 16892
rect 14928 16832 14992 16836
rect 15008 16892 15072 16896
rect 15008 16836 15012 16892
rect 15012 16836 15068 16892
rect 15068 16836 15072 16892
rect 15008 16832 15072 16836
rect 15088 16892 15152 16896
rect 15088 16836 15092 16892
rect 15092 16836 15148 16892
rect 15148 16836 15152 16892
rect 15088 16832 15152 16836
rect 24112 16892 24176 16896
rect 24112 16836 24116 16892
rect 24116 16836 24172 16892
rect 24172 16836 24176 16892
rect 24112 16832 24176 16836
rect 24192 16892 24256 16896
rect 24192 16836 24196 16892
rect 24196 16836 24252 16892
rect 24252 16836 24256 16892
rect 24192 16832 24256 16836
rect 24272 16892 24336 16896
rect 24272 16836 24276 16892
rect 24276 16836 24332 16892
rect 24332 16836 24336 16892
rect 24272 16832 24336 16836
rect 24352 16892 24416 16896
rect 24352 16836 24356 16892
rect 24356 16836 24412 16892
rect 24412 16836 24416 16892
rect 24352 16832 24416 16836
rect 13860 16688 13924 16692
rect 13860 16632 13874 16688
rect 13874 16632 13924 16688
rect 13860 16628 13924 16632
rect 14228 16628 14292 16692
rect 10216 16348 10280 16352
rect 10216 16292 10220 16348
rect 10220 16292 10276 16348
rect 10276 16292 10280 16348
rect 10216 16288 10280 16292
rect 10296 16348 10360 16352
rect 10296 16292 10300 16348
rect 10300 16292 10356 16348
rect 10356 16292 10360 16348
rect 10296 16288 10360 16292
rect 10376 16348 10440 16352
rect 10376 16292 10380 16348
rect 10380 16292 10436 16348
rect 10436 16292 10440 16348
rect 10376 16288 10440 16292
rect 10456 16348 10520 16352
rect 10456 16292 10460 16348
rect 10460 16292 10516 16348
rect 10516 16292 10520 16348
rect 10456 16288 10520 16292
rect 19480 16348 19544 16352
rect 19480 16292 19484 16348
rect 19484 16292 19540 16348
rect 19540 16292 19544 16348
rect 19480 16288 19544 16292
rect 19560 16348 19624 16352
rect 19560 16292 19564 16348
rect 19564 16292 19620 16348
rect 19620 16292 19624 16348
rect 19560 16288 19624 16292
rect 19640 16348 19704 16352
rect 19640 16292 19644 16348
rect 19644 16292 19700 16348
rect 19700 16292 19704 16348
rect 19640 16288 19704 16292
rect 19720 16348 19784 16352
rect 19720 16292 19724 16348
rect 19724 16292 19780 16348
rect 19780 16292 19784 16348
rect 19720 16288 19784 16292
rect 5584 15804 5648 15808
rect 5584 15748 5588 15804
rect 5588 15748 5644 15804
rect 5644 15748 5648 15804
rect 5584 15744 5648 15748
rect 5664 15804 5728 15808
rect 5664 15748 5668 15804
rect 5668 15748 5724 15804
rect 5724 15748 5728 15804
rect 5664 15744 5728 15748
rect 5744 15804 5808 15808
rect 5744 15748 5748 15804
rect 5748 15748 5804 15804
rect 5804 15748 5808 15804
rect 5744 15744 5808 15748
rect 5824 15804 5888 15808
rect 5824 15748 5828 15804
rect 5828 15748 5884 15804
rect 5884 15748 5888 15804
rect 5824 15744 5888 15748
rect 14848 15804 14912 15808
rect 14848 15748 14852 15804
rect 14852 15748 14908 15804
rect 14908 15748 14912 15804
rect 14848 15744 14912 15748
rect 14928 15804 14992 15808
rect 14928 15748 14932 15804
rect 14932 15748 14988 15804
rect 14988 15748 14992 15804
rect 14928 15744 14992 15748
rect 15008 15804 15072 15808
rect 15008 15748 15012 15804
rect 15012 15748 15068 15804
rect 15068 15748 15072 15804
rect 15008 15744 15072 15748
rect 15088 15804 15152 15808
rect 15088 15748 15092 15804
rect 15092 15748 15148 15804
rect 15148 15748 15152 15804
rect 15088 15744 15152 15748
rect 24112 15804 24176 15808
rect 24112 15748 24116 15804
rect 24116 15748 24172 15804
rect 24172 15748 24176 15804
rect 24112 15744 24176 15748
rect 24192 15804 24256 15808
rect 24192 15748 24196 15804
rect 24196 15748 24252 15804
rect 24252 15748 24256 15804
rect 24192 15744 24256 15748
rect 24272 15804 24336 15808
rect 24272 15748 24276 15804
rect 24276 15748 24332 15804
rect 24332 15748 24336 15804
rect 24272 15744 24336 15748
rect 24352 15804 24416 15808
rect 24352 15748 24356 15804
rect 24356 15748 24412 15804
rect 24412 15748 24416 15804
rect 24352 15744 24416 15748
rect 21036 15404 21100 15468
rect 10216 15260 10280 15264
rect 10216 15204 10220 15260
rect 10220 15204 10276 15260
rect 10276 15204 10280 15260
rect 10216 15200 10280 15204
rect 10296 15260 10360 15264
rect 10296 15204 10300 15260
rect 10300 15204 10356 15260
rect 10356 15204 10360 15260
rect 10296 15200 10360 15204
rect 10376 15260 10440 15264
rect 10376 15204 10380 15260
rect 10380 15204 10436 15260
rect 10436 15204 10440 15260
rect 10376 15200 10440 15204
rect 10456 15260 10520 15264
rect 10456 15204 10460 15260
rect 10460 15204 10516 15260
rect 10516 15204 10520 15260
rect 10456 15200 10520 15204
rect 19480 15260 19544 15264
rect 19480 15204 19484 15260
rect 19484 15204 19540 15260
rect 19540 15204 19544 15260
rect 19480 15200 19544 15204
rect 19560 15260 19624 15264
rect 19560 15204 19564 15260
rect 19564 15204 19620 15260
rect 19620 15204 19624 15260
rect 19560 15200 19624 15204
rect 19640 15260 19704 15264
rect 19640 15204 19644 15260
rect 19644 15204 19700 15260
rect 19700 15204 19704 15260
rect 19640 15200 19704 15204
rect 19720 15260 19784 15264
rect 19720 15204 19724 15260
rect 19724 15204 19780 15260
rect 19780 15204 19784 15260
rect 19720 15200 19784 15204
rect 5584 14716 5648 14720
rect 5584 14660 5588 14716
rect 5588 14660 5644 14716
rect 5644 14660 5648 14716
rect 5584 14656 5648 14660
rect 5664 14716 5728 14720
rect 5664 14660 5668 14716
rect 5668 14660 5724 14716
rect 5724 14660 5728 14716
rect 5664 14656 5728 14660
rect 5744 14716 5808 14720
rect 5744 14660 5748 14716
rect 5748 14660 5804 14716
rect 5804 14660 5808 14716
rect 5744 14656 5808 14660
rect 5824 14716 5888 14720
rect 5824 14660 5828 14716
rect 5828 14660 5884 14716
rect 5884 14660 5888 14716
rect 5824 14656 5888 14660
rect 14848 14716 14912 14720
rect 14848 14660 14852 14716
rect 14852 14660 14908 14716
rect 14908 14660 14912 14716
rect 14848 14656 14912 14660
rect 14928 14716 14992 14720
rect 14928 14660 14932 14716
rect 14932 14660 14988 14716
rect 14988 14660 14992 14716
rect 14928 14656 14992 14660
rect 15008 14716 15072 14720
rect 15008 14660 15012 14716
rect 15012 14660 15068 14716
rect 15068 14660 15072 14716
rect 15008 14656 15072 14660
rect 15088 14716 15152 14720
rect 15088 14660 15092 14716
rect 15092 14660 15148 14716
rect 15148 14660 15152 14716
rect 15088 14656 15152 14660
rect 24112 14716 24176 14720
rect 24112 14660 24116 14716
rect 24116 14660 24172 14716
rect 24172 14660 24176 14716
rect 24112 14656 24176 14660
rect 24192 14716 24256 14720
rect 24192 14660 24196 14716
rect 24196 14660 24252 14716
rect 24252 14660 24256 14716
rect 24192 14656 24256 14660
rect 24272 14716 24336 14720
rect 24272 14660 24276 14716
rect 24276 14660 24332 14716
rect 24332 14660 24336 14716
rect 24272 14656 24336 14660
rect 24352 14716 24416 14720
rect 24352 14660 24356 14716
rect 24356 14660 24412 14716
rect 24412 14660 24416 14716
rect 24352 14656 24416 14660
rect 15332 14452 15396 14516
rect 10216 14172 10280 14176
rect 10216 14116 10220 14172
rect 10220 14116 10276 14172
rect 10276 14116 10280 14172
rect 10216 14112 10280 14116
rect 10296 14172 10360 14176
rect 10296 14116 10300 14172
rect 10300 14116 10356 14172
rect 10356 14116 10360 14172
rect 10296 14112 10360 14116
rect 10376 14172 10440 14176
rect 10376 14116 10380 14172
rect 10380 14116 10436 14172
rect 10436 14116 10440 14172
rect 10376 14112 10440 14116
rect 10456 14172 10520 14176
rect 10456 14116 10460 14172
rect 10460 14116 10516 14172
rect 10516 14116 10520 14172
rect 10456 14112 10520 14116
rect 19480 14172 19544 14176
rect 19480 14116 19484 14172
rect 19484 14116 19540 14172
rect 19540 14116 19544 14172
rect 19480 14112 19544 14116
rect 19560 14172 19624 14176
rect 19560 14116 19564 14172
rect 19564 14116 19620 14172
rect 19620 14116 19624 14172
rect 19560 14112 19624 14116
rect 19640 14172 19704 14176
rect 19640 14116 19644 14172
rect 19644 14116 19700 14172
rect 19700 14116 19704 14172
rect 19640 14112 19704 14116
rect 19720 14172 19784 14176
rect 19720 14116 19724 14172
rect 19724 14116 19780 14172
rect 19780 14116 19784 14172
rect 19720 14112 19784 14116
rect 5584 13628 5648 13632
rect 5584 13572 5588 13628
rect 5588 13572 5644 13628
rect 5644 13572 5648 13628
rect 5584 13568 5648 13572
rect 5664 13628 5728 13632
rect 5664 13572 5668 13628
rect 5668 13572 5724 13628
rect 5724 13572 5728 13628
rect 5664 13568 5728 13572
rect 5744 13628 5808 13632
rect 5744 13572 5748 13628
rect 5748 13572 5804 13628
rect 5804 13572 5808 13628
rect 5744 13568 5808 13572
rect 5824 13628 5888 13632
rect 5824 13572 5828 13628
rect 5828 13572 5884 13628
rect 5884 13572 5888 13628
rect 5824 13568 5888 13572
rect 14848 13628 14912 13632
rect 14848 13572 14852 13628
rect 14852 13572 14908 13628
rect 14908 13572 14912 13628
rect 14848 13568 14912 13572
rect 14928 13628 14992 13632
rect 14928 13572 14932 13628
rect 14932 13572 14988 13628
rect 14988 13572 14992 13628
rect 14928 13568 14992 13572
rect 15008 13628 15072 13632
rect 15008 13572 15012 13628
rect 15012 13572 15068 13628
rect 15068 13572 15072 13628
rect 15008 13568 15072 13572
rect 15088 13628 15152 13632
rect 15088 13572 15092 13628
rect 15092 13572 15148 13628
rect 15148 13572 15152 13628
rect 15088 13568 15152 13572
rect 24112 13628 24176 13632
rect 24112 13572 24116 13628
rect 24116 13572 24172 13628
rect 24172 13572 24176 13628
rect 24112 13568 24176 13572
rect 24192 13628 24256 13632
rect 24192 13572 24196 13628
rect 24196 13572 24252 13628
rect 24252 13572 24256 13628
rect 24192 13568 24256 13572
rect 24272 13628 24336 13632
rect 24272 13572 24276 13628
rect 24276 13572 24332 13628
rect 24332 13572 24336 13628
rect 24272 13568 24336 13572
rect 24352 13628 24416 13632
rect 24352 13572 24356 13628
rect 24356 13572 24412 13628
rect 24412 13572 24416 13628
rect 24352 13568 24416 13572
rect 15332 13228 15396 13292
rect 10216 13084 10280 13088
rect 10216 13028 10220 13084
rect 10220 13028 10276 13084
rect 10276 13028 10280 13084
rect 10216 13024 10280 13028
rect 10296 13084 10360 13088
rect 10296 13028 10300 13084
rect 10300 13028 10356 13084
rect 10356 13028 10360 13084
rect 10296 13024 10360 13028
rect 10376 13084 10440 13088
rect 10376 13028 10380 13084
rect 10380 13028 10436 13084
rect 10436 13028 10440 13084
rect 10376 13024 10440 13028
rect 10456 13084 10520 13088
rect 10456 13028 10460 13084
rect 10460 13028 10516 13084
rect 10516 13028 10520 13084
rect 10456 13024 10520 13028
rect 19480 13084 19544 13088
rect 19480 13028 19484 13084
rect 19484 13028 19540 13084
rect 19540 13028 19544 13084
rect 19480 13024 19544 13028
rect 19560 13084 19624 13088
rect 19560 13028 19564 13084
rect 19564 13028 19620 13084
rect 19620 13028 19624 13084
rect 19560 13024 19624 13028
rect 19640 13084 19704 13088
rect 19640 13028 19644 13084
rect 19644 13028 19700 13084
rect 19700 13028 19704 13084
rect 19640 13024 19704 13028
rect 19720 13084 19784 13088
rect 19720 13028 19724 13084
rect 19724 13028 19780 13084
rect 19780 13028 19784 13084
rect 19720 13024 19784 13028
rect 5584 12540 5648 12544
rect 5584 12484 5588 12540
rect 5588 12484 5644 12540
rect 5644 12484 5648 12540
rect 5584 12480 5648 12484
rect 5664 12540 5728 12544
rect 5664 12484 5668 12540
rect 5668 12484 5724 12540
rect 5724 12484 5728 12540
rect 5664 12480 5728 12484
rect 5744 12540 5808 12544
rect 5744 12484 5748 12540
rect 5748 12484 5804 12540
rect 5804 12484 5808 12540
rect 5744 12480 5808 12484
rect 5824 12540 5888 12544
rect 5824 12484 5828 12540
rect 5828 12484 5884 12540
rect 5884 12484 5888 12540
rect 5824 12480 5888 12484
rect 14848 12540 14912 12544
rect 14848 12484 14852 12540
rect 14852 12484 14908 12540
rect 14908 12484 14912 12540
rect 14848 12480 14912 12484
rect 14928 12540 14992 12544
rect 14928 12484 14932 12540
rect 14932 12484 14988 12540
rect 14988 12484 14992 12540
rect 14928 12480 14992 12484
rect 15008 12540 15072 12544
rect 15008 12484 15012 12540
rect 15012 12484 15068 12540
rect 15068 12484 15072 12540
rect 15008 12480 15072 12484
rect 15088 12540 15152 12544
rect 15088 12484 15092 12540
rect 15092 12484 15148 12540
rect 15148 12484 15152 12540
rect 15088 12480 15152 12484
rect 24112 12540 24176 12544
rect 24112 12484 24116 12540
rect 24116 12484 24172 12540
rect 24172 12484 24176 12540
rect 24112 12480 24176 12484
rect 24192 12540 24256 12544
rect 24192 12484 24196 12540
rect 24196 12484 24252 12540
rect 24252 12484 24256 12540
rect 24192 12480 24256 12484
rect 24272 12540 24336 12544
rect 24272 12484 24276 12540
rect 24276 12484 24332 12540
rect 24332 12484 24336 12540
rect 24272 12480 24336 12484
rect 24352 12540 24416 12544
rect 24352 12484 24356 12540
rect 24356 12484 24412 12540
rect 24412 12484 24416 12540
rect 24352 12480 24416 12484
rect 17540 12064 17604 12068
rect 17540 12008 17554 12064
rect 17554 12008 17604 12064
rect 17540 12004 17604 12008
rect 10216 11996 10280 12000
rect 10216 11940 10220 11996
rect 10220 11940 10276 11996
rect 10276 11940 10280 11996
rect 10216 11936 10280 11940
rect 10296 11996 10360 12000
rect 10296 11940 10300 11996
rect 10300 11940 10356 11996
rect 10356 11940 10360 11996
rect 10296 11936 10360 11940
rect 10376 11996 10440 12000
rect 10376 11940 10380 11996
rect 10380 11940 10436 11996
rect 10436 11940 10440 11996
rect 10376 11936 10440 11940
rect 10456 11996 10520 12000
rect 10456 11940 10460 11996
rect 10460 11940 10516 11996
rect 10516 11940 10520 11996
rect 10456 11936 10520 11940
rect 19480 11996 19544 12000
rect 19480 11940 19484 11996
rect 19484 11940 19540 11996
rect 19540 11940 19544 11996
rect 19480 11936 19544 11940
rect 19560 11996 19624 12000
rect 19560 11940 19564 11996
rect 19564 11940 19620 11996
rect 19620 11940 19624 11996
rect 19560 11936 19624 11940
rect 19640 11996 19704 12000
rect 19640 11940 19644 11996
rect 19644 11940 19700 11996
rect 19700 11940 19704 11996
rect 19640 11936 19704 11940
rect 19720 11996 19784 12000
rect 19720 11940 19724 11996
rect 19724 11940 19780 11996
rect 19780 11940 19784 11996
rect 19720 11936 19784 11940
rect 5584 11452 5648 11456
rect 5584 11396 5588 11452
rect 5588 11396 5644 11452
rect 5644 11396 5648 11452
rect 5584 11392 5648 11396
rect 5664 11452 5728 11456
rect 5664 11396 5668 11452
rect 5668 11396 5724 11452
rect 5724 11396 5728 11452
rect 5664 11392 5728 11396
rect 5744 11452 5808 11456
rect 5744 11396 5748 11452
rect 5748 11396 5804 11452
rect 5804 11396 5808 11452
rect 5744 11392 5808 11396
rect 5824 11452 5888 11456
rect 5824 11396 5828 11452
rect 5828 11396 5884 11452
rect 5884 11396 5888 11452
rect 5824 11392 5888 11396
rect 14848 11452 14912 11456
rect 14848 11396 14852 11452
rect 14852 11396 14908 11452
rect 14908 11396 14912 11452
rect 14848 11392 14912 11396
rect 14928 11452 14992 11456
rect 14928 11396 14932 11452
rect 14932 11396 14988 11452
rect 14988 11396 14992 11452
rect 14928 11392 14992 11396
rect 15008 11452 15072 11456
rect 15008 11396 15012 11452
rect 15012 11396 15068 11452
rect 15068 11396 15072 11452
rect 15008 11392 15072 11396
rect 15088 11452 15152 11456
rect 15088 11396 15092 11452
rect 15092 11396 15148 11452
rect 15148 11396 15152 11452
rect 15088 11392 15152 11396
rect 24112 11452 24176 11456
rect 24112 11396 24116 11452
rect 24116 11396 24172 11452
rect 24172 11396 24176 11452
rect 24112 11392 24176 11396
rect 24192 11452 24256 11456
rect 24192 11396 24196 11452
rect 24196 11396 24252 11452
rect 24252 11396 24256 11452
rect 24192 11392 24256 11396
rect 24272 11452 24336 11456
rect 24272 11396 24276 11452
rect 24276 11396 24332 11452
rect 24332 11396 24336 11452
rect 24272 11392 24336 11396
rect 24352 11452 24416 11456
rect 24352 11396 24356 11452
rect 24356 11396 24412 11452
rect 24412 11396 24416 11452
rect 24352 11392 24416 11396
rect 11100 11112 11164 11116
rect 11100 11056 11150 11112
rect 11150 11056 11164 11112
rect 11100 11052 11164 11056
rect 10216 10908 10280 10912
rect 10216 10852 10220 10908
rect 10220 10852 10276 10908
rect 10276 10852 10280 10908
rect 10216 10848 10280 10852
rect 10296 10908 10360 10912
rect 10296 10852 10300 10908
rect 10300 10852 10356 10908
rect 10356 10852 10360 10908
rect 10296 10848 10360 10852
rect 10376 10908 10440 10912
rect 10376 10852 10380 10908
rect 10380 10852 10436 10908
rect 10436 10852 10440 10908
rect 10376 10848 10440 10852
rect 10456 10908 10520 10912
rect 10456 10852 10460 10908
rect 10460 10852 10516 10908
rect 10516 10852 10520 10908
rect 10456 10848 10520 10852
rect 19480 10908 19544 10912
rect 19480 10852 19484 10908
rect 19484 10852 19540 10908
rect 19540 10852 19544 10908
rect 19480 10848 19544 10852
rect 19560 10908 19624 10912
rect 19560 10852 19564 10908
rect 19564 10852 19620 10908
rect 19620 10852 19624 10908
rect 19560 10848 19624 10852
rect 19640 10908 19704 10912
rect 19640 10852 19644 10908
rect 19644 10852 19700 10908
rect 19700 10852 19704 10908
rect 19640 10848 19704 10852
rect 19720 10908 19784 10912
rect 19720 10852 19724 10908
rect 19724 10852 19780 10908
rect 19780 10852 19784 10908
rect 19720 10848 19784 10852
rect 5584 10364 5648 10368
rect 5584 10308 5588 10364
rect 5588 10308 5644 10364
rect 5644 10308 5648 10364
rect 5584 10304 5648 10308
rect 5664 10364 5728 10368
rect 5664 10308 5668 10364
rect 5668 10308 5724 10364
rect 5724 10308 5728 10364
rect 5664 10304 5728 10308
rect 5744 10364 5808 10368
rect 5744 10308 5748 10364
rect 5748 10308 5804 10364
rect 5804 10308 5808 10364
rect 5744 10304 5808 10308
rect 5824 10364 5888 10368
rect 5824 10308 5828 10364
rect 5828 10308 5884 10364
rect 5884 10308 5888 10364
rect 5824 10304 5888 10308
rect 14848 10364 14912 10368
rect 14848 10308 14852 10364
rect 14852 10308 14908 10364
rect 14908 10308 14912 10364
rect 14848 10304 14912 10308
rect 14928 10364 14992 10368
rect 14928 10308 14932 10364
rect 14932 10308 14988 10364
rect 14988 10308 14992 10364
rect 14928 10304 14992 10308
rect 15008 10364 15072 10368
rect 15008 10308 15012 10364
rect 15012 10308 15068 10364
rect 15068 10308 15072 10364
rect 15008 10304 15072 10308
rect 15088 10364 15152 10368
rect 15088 10308 15092 10364
rect 15092 10308 15148 10364
rect 15148 10308 15152 10364
rect 15088 10304 15152 10308
rect 24112 10364 24176 10368
rect 24112 10308 24116 10364
rect 24116 10308 24172 10364
rect 24172 10308 24176 10364
rect 24112 10304 24176 10308
rect 24192 10364 24256 10368
rect 24192 10308 24196 10364
rect 24196 10308 24252 10364
rect 24252 10308 24256 10364
rect 24192 10304 24256 10308
rect 24272 10364 24336 10368
rect 24272 10308 24276 10364
rect 24276 10308 24332 10364
rect 24332 10308 24336 10364
rect 24272 10304 24336 10308
rect 24352 10364 24416 10368
rect 24352 10308 24356 10364
rect 24356 10308 24412 10364
rect 24412 10308 24416 10364
rect 24352 10304 24416 10308
rect 10216 9820 10280 9824
rect 10216 9764 10220 9820
rect 10220 9764 10276 9820
rect 10276 9764 10280 9820
rect 10216 9760 10280 9764
rect 10296 9820 10360 9824
rect 10296 9764 10300 9820
rect 10300 9764 10356 9820
rect 10356 9764 10360 9820
rect 10296 9760 10360 9764
rect 10376 9820 10440 9824
rect 10376 9764 10380 9820
rect 10380 9764 10436 9820
rect 10436 9764 10440 9820
rect 10376 9760 10440 9764
rect 10456 9820 10520 9824
rect 10456 9764 10460 9820
rect 10460 9764 10516 9820
rect 10516 9764 10520 9820
rect 10456 9760 10520 9764
rect 19480 9820 19544 9824
rect 19480 9764 19484 9820
rect 19484 9764 19540 9820
rect 19540 9764 19544 9820
rect 19480 9760 19544 9764
rect 19560 9820 19624 9824
rect 19560 9764 19564 9820
rect 19564 9764 19620 9820
rect 19620 9764 19624 9820
rect 19560 9760 19624 9764
rect 19640 9820 19704 9824
rect 19640 9764 19644 9820
rect 19644 9764 19700 9820
rect 19700 9764 19704 9820
rect 19640 9760 19704 9764
rect 19720 9820 19784 9824
rect 19720 9764 19724 9820
rect 19724 9764 19780 9820
rect 19780 9764 19784 9820
rect 19720 9760 19784 9764
rect 5584 9276 5648 9280
rect 5584 9220 5588 9276
rect 5588 9220 5644 9276
rect 5644 9220 5648 9276
rect 5584 9216 5648 9220
rect 5664 9276 5728 9280
rect 5664 9220 5668 9276
rect 5668 9220 5724 9276
rect 5724 9220 5728 9276
rect 5664 9216 5728 9220
rect 5744 9276 5808 9280
rect 5744 9220 5748 9276
rect 5748 9220 5804 9276
rect 5804 9220 5808 9276
rect 5744 9216 5808 9220
rect 5824 9276 5888 9280
rect 5824 9220 5828 9276
rect 5828 9220 5884 9276
rect 5884 9220 5888 9276
rect 5824 9216 5888 9220
rect 14848 9276 14912 9280
rect 14848 9220 14852 9276
rect 14852 9220 14908 9276
rect 14908 9220 14912 9276
rect 14848 9216 14912 9220
rect 14928 9276 14992 9280
rect 14928 9220 14932 9276
rect 14932 9220 14988 9276
rect 14988 9220 14992 9276
rect 14928 9216 14992 9220
rect 15008 9276 15072 9280
rect 15008 9220 15012 9276
rect 15012 9220 15068 9276
rect 15068 9220 15072 9276
rect 15008 9216 15072 9220
rect 15088 9276 15152 9280
rect 15088 9220 15092 9276
rect 15092 9220 15148 9276
rect 15148 9220 15152 9276
rect 15088 9216 15152 9220
rect 24112 9276 24176 9280
rect 24112 9220 24116 9276
rect 24116 9220 24172 9276
rect 24172 9220 24176 9276
rect 24112 9216 24176 9220
rect 24192 9276 24256 9280
rect 24192 9220 24196 9276
rect 24196 9220 24252 9276
rect 24252 9220 24256 9276
rect 24192 9216 24256 9220
rect 24272 9276 24336 9280
rect 24272 9220 24276 9276
rect 24276 9220 24332 9276
rect 24332 9220 24336 9276
rect 24272 9216 24336 9220
rect 24352 9276 24416 9280
rect 24352 9220 24356 9276
rect 24356 9220 24412 9276
rect 24412 9220 24416 9276
rect 24352 9216 24416 9220
rect 10216 8732 10280 8736
rect 10216 8676 10220 8732
rect 10220 8676 10276 8732
rect 10276 8676 10280 8732
rect 10216 8672 10280 8676
rect 10296 8732 10360 8736
rect 10296 8676 10300 8732
rect 10300 8676 10356 8732
rect 10356 8676 10360 8732
rect 10296 8672 10360 8676
rect 10376 8732 10440 8736
rect 10376 8676 10380 8732
rect 10380 8676 10436 8732
rect 10436 8676 10440 8732
rect 10376 8672 10440 8676
rect 10456 8732 10520 8736
rect 10456 8676 10460 8732
rect 10460 8676 10516 8732
rect 10516 8676 10520 8732
rect 10456 8672 10520 8676
rect 19480 8732 19544 8736
rect 19480 8676 19484 8732
rect 19484 8676 19540 8732
rect 19540 8676 19544 8732
rect 19480 8672 19544 8676
rect 19560 8732 19624 8736
rect 19560 8676 19564 8732
rect 19564 8676 19620 8732
rect 19620 8676 19624 8732
rect 19560 8672 19624 8676
rect 19640 8732 19704 8736
rect 19640 8676 19644 8732
rect 19644 8676 19700 8732
rect 19700 8676 19704 8732
rect 19640 8672 19704 8676
rect 19720 8732 19784 8736
rect 19720 8676 19724 8732
rect 19724 8676 19780 8732
rect 19780 8676 19784 8732
rect 19720 8672 19784 8676
rect 5584 8188 5648 8192
rect 5584 8132 5588 8188
rect 5588 8132 5644 8188
rect 5644 8132 5648 8188
rect 5584 8128 5648 8132
rect 5664 8188 5728 8192
rect 5664 8132 5668 8188
rect 5668 8132 5724 8188
rect 5724 8132 5728 8188
rect 5664 8128 5728 8132
rect 5744 8188 5808 8192
rect 5744 8132 5748 8188
rect 5748 8132 5804 8188
rect 5804 8132 5808 8188
rect 5744 8128 5808 8132
rect 5824 8188 5888 8192
rect 5824 8132 5828 8188
rect 5828 8132 5884 8188
rect 5884 8132 5888 8188
rect 5824 8128 5888 8132
rect 14848 8188 14912 8192
rect 14848 8132 14852 8188
rect 14852 8132 14908 8188
rect 14908 8132 14912 8188
rect 14848 8128 14912 8132
rect 14928 8188 14992 8192
rect 14928 8132 14932 8188
rect 14932 8132 14988 8188
rect 14988 8132 14992 8188
rect 14928 8128 14992 8132
rect 15008 8188 15072 8192
rect 15008 8132 15012 8188
rect 15012 8132 15068 8188
rect 15068 8132 15072 8188
rect 15008 8128 15072 8132
rect 15088 8188 15152 8192
rect 15088 8132 15092 8188
rect 15092 8132 15148 8188
rect 15148 8132 15152 8188
rect 15088 8128 15152 8132
rect 24112 8188 24176 8192
rect 24112 8132 24116 8188
rect 24116 8132 24172 8188
rect 24172 8132 24176 8188
rect 24112 8128 24176 8132
rect 24192 8188 24256 8192
rect 24192 8132 24196 8188
rect 24196 8132 24252 8188
rect 24252 8132 24256 8188
rect 24192 8128 24256 8132
rect 24272 8188 24336 8192
rect 24272 8132 24276 8188
rect 24276 8132 24332 8188
rect 24332 8132 24336 8188
rect 24272 8128 24336 8132
rect 24352 8188 24416 8192
rect 24352 8132 24356 8188
rect 24356 8132 24412 8188
rect 24412 8132 24416 8188
rect 24352 8128 24416 8132
rect 11100 7924 11164 7988
rect 10216 7644 10280 7648
rect 10216 7588 10220 7644
rect 10220 7588 10276 7644
rect 10276 7588 10280 7644
rect 10216 7584 10280 7588
rect 10296 7644 10360 7648
rect 10296 7588 10300 7644
rect 10300 7588 10356 7644
rect 10356 7588 10360 7644
rect 10296 7584 10360 7588
rect 10376 7644 10440 7648
rect 10376 7588 10380 7644
rect 10380 7588 10436 7644
rect 10436 7588 10440 7644
rect 10376 7584 10440 7588
rect 10456 7644 10520 7648
rect 10456 7588 10460 7644
rect 10460 7588 10516 7644
rect 10516 7588 10520 7644
rect 10456 7584 10520 7588
rect 19480 7644 19544 7648
rect 19480 7588 19484 7644
rect 19484 7588 19540 7644
rect 19540 7588 19544 7644
rect 19480 7584 19544 7588
rect 19560 7644 19624 7648
rect 19560 7588 19564 7644
rect 19564 7588 19620 7644
rect 19620 7588 19624 7644
rect 19560 7584 19624 7588
rect 19640 7644 19704 7648
rect 19640 7588 19644 7644
rect 19644 7588 19700 7644
rect 19700 7588 19704 7644
rect 19640 7584 19704 7588
rect 19720 7644 19784 7648
rect 19720 7588 19724 7644
rect 19724 7588 19780 7644
rect 19780 7588 19784 7644
rect 19720 7584 19784 7588
rect 5584 7100 5648 7104
rect 5584 7044 5588 7100
rect 5588 7044 5644 7100
rect 5644 7044 5648 7100
rect 5584 7040 5648 7044
rect 5664 7100 5728 7104
rect 5664 7044 5668 7100
rect 5668 7044 5724 7100
rect 5724 7044 5728 7100
rect 5664 7040 5728 7044
rect 5744 7100 5808 7104
rect 5744 7044 5748 7100
rect 5748 7044 5804 7100
rect 5804 7044 5808 7100
rect 5744 7040 5808 7044
rect 5824 7100 5888 7104
rect 5824 7044 5828 7100
rect 5828 7044 5884 7100
rect 5884 7044 5888 7100
rect 5824 7040 5888 7044
rect 14848 7100 14912 7104
rect 14848 7044 14852 7100
rect 14852 7044 14908 7100
rect 14908 7044 14912 7100
rect 14848 7040 14912 7044
rect 14928 7100 14992 7104
rect 14928 7044 14932 7100
rect 14932 7044 14988 7100
rect 14988 7044 14992 7100
rect 14928 7040 14992 7044
rect 15008 7100 15072 7104
rect 15008 7044 15012 7100
rect 15012 7044 15068 7100
rect 15068 7044 15072 7100
rect 15008 7040 15072 7044
rect 15088 7100 15152 7104
rect 15088 7044 15092 7100
rect 15092 7044 15148 7100
rect 15148 7044 15152 7100
rect 15088 7040 15152 7044
rect 24112 7100 24176 7104
rect 24112 7044 24116 7100
rect 24116 7044 24172 7100
rect 24172 7044 24176 7100
rect 24112 7040 24176 7044
rect 24192 7100 24256 7104
rect 24192 7044 24196 7100
rect 24196 7044 24252 7100
rect 24252 7044 24256 7100
rect 24192 7040 24256 7044
rect 24272 7100 24336 7104
rect 24272 7044 24276 7100
rect 24276 7044 24332 7100
rect 24332 7044 24336 7100
rect 24272 7040 24336 7044
rect 24352 7100 24416 7104
rect 24352 7044 24356 7100
rect 24356 7044 24412 7100
rect 24412 7044 24416 7100
rect 24352 7040 24416 7044
rect 10216 6556 10280 6560
rect 10216 6500 10220 6556
rect 10220 6500 10276 6556
rect 10276 6500 10280 6556
rect 10216 6496 10280 6500
rect 10296 6556 10360 6560
rect 10296 6500 10300 6556
rect 10300 6500 10356 6556
rect 10356 6500 10360 6556
rect 10296 6496 10360 6500
rect 10376 6556 10440 6560
rect 10376 6500 10380 6556
rect 10380 6500 10436 6556
rect 10436 6500 10440 6556
rect 10376 6496 10440 6500
rect 10456 6556 10520 6560
rect 10456 6500 10460 6556
rect 10460 6500 10516 6556
rect 10516 6500 10520 6556
rect 10456 6496 10520 6500
rect 19480 6556 19544 6560
rect 19480 6500 19484 6556
rect 19484 6500 19540 6556
rect 19540 6500 19544 6556
rect 19480 6496 19544 6500
rect 19560 6556 19624 6560
rect 19560 6500 19564 6556
rect 19564 6500 19620 6556
rect 19620 6500 19624 6556
rect 19560 6496 19624 6500
rect 19640 6556 19704 6560
rect 19640 6500 19644 6556
rect 19644 6500 19700 6556
rect 19700 6500 19704 6556
rect 19640 6496 19704 6500
rect 19720 6556 19784 6560
rect 19720 6500 19724 6556
rect 19724 6500 19780 6556
rect 19780 6500 19784 6556
rect 19720 6496 19784 6500
rect 5584 6012 5648 6016
rect 5584 5956 5588 6012
rect 5588 5956 5644 6012
rect 5644 5956 5648 6012
rect 5584 5952 5648 5956
rect 5664 6012 5728 6016
rect 5664 5956 5668 6012
rect 5668 5956 5724 6012
rect 5724 5956 5728 6012
rect 5664 5952 5728 5956
rect 5744 6012 5808 6016
rect 5744 5956 5748 6012
rect 5748 5956 5804 6012
rect 5804 5956 5808 6012
rect 5744 5952 5808 5956
rect 5824 6012 5888 6016
rect 5824 5956 5828 6012
rect 5828 5956 5884 6012
rect 5884 5956 5888 6012
rect 5824 5952 5888 5956
rect 14848 6012 14912 6016
rect 14848 5956 14852 6012
rect 14852 5956 14908 6012
rect 14908 5956 14912 6012
rect 14848 5952 14912 5956
rect 14928 6012 14992 6016
rect 14928 5956 14932 6012
rect 14932 5956 14988 6012
rect 14988 5956 14992 6012
rect 14928 5952 14992 5956
rect 15008 6012 15072 6016
rect 15008 5956 15012 6012
rect 15012 5956 15068 6012
rect 15068 5956 15072 6012
rect 15008 5952 15072 5956
rect 15088 6012 15152 6016
rect 15088 5956 15092 6012
rect 15092 5956 15148 6012
rect 15148 5956 15152 6012
rect 15088 5952 15152 5956
rect 24112 6012 24176 6016
rect 24112 5956 24116 6012
rect 24116 5956 24172 6012
rect 24172 5956 24176 6012
rect 24112 5952 24176 5956
rect 24192 6012 24256 6016
rect 24192 5956 24196 6012
rect 24196 5956 24252 6012
rect 24252 5956 24256 6012
rect 24192 5952 24256 5956
rect 24272 6012 24336 6016
rect 24272 5956 24276 6012
rect 24276 5956 24332 6012
rect 24332 5956 24336 6012
rect 24272 5952 24336 5956
rect 24352 6012 24416 6016
rect 24352 5956 24356 6012
rect 24356 5956 24412 6012
rect 24412 5956 24416 6012
rect 24352 5952 24416 5956
rect 14228 5884 14292 5948
rect 10216 5468 10280 5472
rect 10216 5412 10220 5468
rect 10220 5412 10276 5468
rect 10276 5412 10280 5468
rect 10216 5408 10280 5412
rect 10296 5468 10360 5472
rect 10296 5412 10300 5468
rect 10300 5412 10356 5468
rect 10356 5412 10360 5468
rect 10296 5408 10360 5412
rect 10376 5468 10440 5472
rect 10376 5412 10380 5468
rect 10380 5412 10436 5468
rect 10436 5412 10440 5468
rect 10376 5408 10440 5412
rect 10456 5468 10520 5472
rect 10456 5412 10460 5468
rect 10460 5412 10516 5468
rect 10516 5412 10520 5468
rect 10456 5408 10520 5412
rect 19480 5468 19544 5472
rect 19480 5412 19484 5468
rect 19484 5412 19540 5468
rect 19540 5412 19544 5468
rect 19480 5408 19544 5412
rect 19560 5468 19624 5472
rect 19560 5412 19564 5468
rect 19564 5412 19620 5468
rect 19620 5412 19624 5468
rect 19560 5408 19624 5412
rect 19640 5468 19704 5472
rect 19640 5412 19644 5468
rect 19644 5412 19700 5468
rect 19700 5412 19704 5468
rect 19640 5408 19704 5412
rect 19720 5468 19784 5472
rect 19720 5412 19724 5468
rect 19724 5412 19780 5468
rect 19780 5412 19784 5468
rect 19720 5408 19784 5412
rect 5584 4924 5648 4928
rect 5584 4868 5588 4924
rect 5588 4868 5644 4924
rect 5644 4868 5648 4924
rect 5584 4864 5648 4868
rect 5664 4924 5728 4928
rect 5664 4868 5668 4924
rect 5668 4868 5724 4924
rect 5724 4868 5728 4924
rect 5664 4864 5728 4868
rect 5744 4924 5808 4928
rect 5744 4868 5748 4924
rect 5748 4868 5804 4924
rect 5804 4868 5808 4924
rect 5744 4864 5808 4868
rect 5824 4924 5888 4928
rect 5824 4868 5828 4924
rect 5828 4868 5884 4924
rect 5884 4868 5888 4924
rect 5824 4864 5888 4868
rect 14848 4924 14912 4928
rect 14848 4868 14852 4924
rect 14852 4868 14908 4924
rect 14908 4868 14912 4924
rect 14848 4864 14912 4868
rect 14928 4924 14992 4928
rect 14928 4868 14932 4924
rect 14932 4868 14988 4924
rect 14988 4868 14992 4924
rect 14928 4864 14992 4868
rect 15008 4924 15072 4928
rect 15008 4868 15012 4924
rect 15012 4868 15068 4924
rect 15068 4868 15072 4924
rect 15008 4864 15072 4868
rect 15088 4924 15152 4928
rect 15088 4868 15092 4924
rect 15092 4868 15148 4924
rect 15148 4868 15152 4924
rect 15088 4864 15152 4868
rect 24112 4924 24176 4928
rect 24112 4868 24116 4924
rect 24116 4868 24172 4924
rect 24172 4868 24176 4924
rect 24112 4864 24176 4868
rect 24192 4924 24256 4928
rect 24192 4868 24196 4924
rect 24196 4868 24252 4924
rect 24252 4868 24256 4924
rect 24192 4864 24256 4868
rect 24272 4924 24336 4928
rect 24272 4868 24276 4924
rect 24276 4868 24332 4924
rect 24332 4868 24336 4924
rect 24272 4864 24336 4868
rect 24352 4924 24416 4928
rect 24352 4868 24356 4924
rect 24356 4868 24412 4924
rect 24412 4868 24416 4924
rect 24352 4864 24416 4868
rect 10216 4380 10280 4384
rect 10216 4324 10220 4380
rect 10220 4324 10276 4380
rect 10276 4324 10280 4380
rect 10216 4320 10280 4324
rect 10296 4380 10360 4384
rect 10296 4324 10300 4380
rect 10300 4324 10356 4380
rect 10356 4324 10360 4380
rect 10296 4320 10360 4324
rect 10376 4380 10440 4384
rect 10376 4324 10380 4380
rect 10380 4324 10436 4380
rect 10436 4324 10440 4380
rect 10376 4320 10440 4324
rect 10456 4380 10520 4384
rect 10456 4324 10460 4380
rect 10460 4324 10516 4380
rect 10516 4324 10520 4380
rect 10456 4320 10520 4324
rect 19480 4380 19544 4384
rect 19480 4324 19484 4380
rect 19484 4324 19540 4380
rect 19540 4324 19544 4380
rect 19480 4320 19544 4324
rect 19560 4380 19624 4384
rect 19560 4324 19564 4380
rect 19564 4324 19620 4380
rect 19620 4324 19624 4380
rect 19560 4320 19624 4324
rect 19640 4380 19704 4384
rect 19640 4324 19644 4380
rect 19644 4324 19700 4380
rect 19700 4324 19704 4380
rect 19640 4320 19704 4324
rect 19720 4380 19784 4384
rect 19720 4324 19724 4380
rect 19724 4324 19780 4380
rect 19780 4324 19784 4380
rect 19720 4320 19784 4324
rect 5584 3836 5648 3840
rect 5584 3780 5588 3836
rect 5588 3780 5644 3836
rect 5644 3780 5648 3836
rect 5584 3776 5648 3780
rect 5664 3836 5728 3840
rect 5664 3780 5668 3836
rect 5668 3780 5724 3836
rect 5724 3780 5728 3836
rect 5664 3776 5728 3780
rect 5744 3836 5808 3840
rect 5744 3780 5748 3836
rect 5748 3780 5804 3836
rect 5804 3780 5808 3836
rect 5744 3776 5808 3780
rect 5824 3836 5888 3840
rect 5824 3780 5828 3836
rect 5828 3780 5884 3836
rect 5884 3780 5888 3836
rect 5824 3776 5888 3780
rect 14848 3836 14912 3840
rect 14848 3780 14852 3836
rect 14852 3780 14908 3836
rect 14908 3780 14912 3836
rect 14848 3776 14912 3780
rect 14928 3836 14992 3840
rect 14928 3780 14932 3836
rect 14932 3780 14988 3836
rect 14988 3780 14992 3836
rect 14928 3776 14992 3780
rect 15008 3836 15072 3840
rect 15008 3780 15012 3836
rect 15012 3780 15068 3836
rect 15068 3780 15072 3836
rect 15008 3776 15072 3780
rect 15088 3836 15152 3840
rect 15088 3780 15092 3836
rect 15092 3780 15148 3836
rect 15148 3780 15152 3836
rect 15088 3776 15152 3780
rect 24112 3836 24176 3840
rect 24112 3780 24116 3836
rect 24116 3780 24172 3836
rect 24172 3780 24176 3836
rect 24112 3776 24176 3780
rect 24192 3836 24256 3840
rect 24192 3780 24196 3836
rect 24196 3780 24252 3836
rect 24252 3780 24256 3836
rect 24192 3776 24256 3780
rect 24272 3836 24336 3840
rect 24272 3780 24276 3836
rect 24276 3780 24332 3836
rect 24332 3780 24336 3836
rect 24272 3776 24336 3780
rect 24352 3836 24416 3840
rect 24352 3780 24356 3836
rect 24356 3780 24412 3836
rect 24412 3780 24416 3836
rect 24352 3776 24416 3780
rect 13860 3436 13924 3500
rect 10216 3292 10280 3296
rect 10216 3236 10220 3292
rect 10220 3236 10276 3292
rect 10276 3236 10280 3292
rect 10216 3232 10280 3236
rect 10296 3292 10360 3296
rect 10296 3236 10300 3292
rect 10300 3236 10356 3292
rect 10356 3236 10360 3292
rect 10296 3232 10360 3236
rect 10376 3292 10440 3296
rect 10376 3236 10380 3292
rect 10380 3236 10436 3292
rect 10436 3236 10440 3292
rect 10376 3232 10440 3236
rect 10456 3292 10520 3296
rect 10456 3236 10460 3292
rect 10460 3236 10516 3292
rect 10516 3236 10520 3292
rect 10456 3232 10520 3236
rect 19480 3292 19544 3296
rect 19480 3236 19484 3292
rect 19484 3236 19540 3292
rect 19540 3236 19544 3292
rect 19480 3232 19544 3236
rect 19560 3292 19624 3296
rect 19560 3236 19564 3292
rect 19564 3236 19620 3292
rect 19620 3236 19624 3292
rect 19560 3232 19624 3236
rect 19640 3292 19704 3296
rect 19640 3236 19644 3292
rect 19644 3236 19700 3292
rect 19700 3236 19704 3292
rect 19640 3232 19704 3236
rect 19720 3292 19784 3296
rect 19720 3236 19724 3292
rect 19724 3236 19780 3292
rect 19780 3236 19784 3292
rect 19720 3232 19784 3236
rect 5584 2748 5648 2752
rect 5584 2692 5588 2748
rect 5588 2692 5644 2748
rect 5644 2692 5648 2748
rect 5584 2688 5648 2692
rect 5664 2748 5728 2752
rect 5664 2692 5668 2748
rect 5668 2692 5724 2748
rect 5724 2692 5728 2748
rect 5664 2688 5728 2692
rect 5744 2748 5808 2752
rect 5744 2692 5748 2748
rect 5748 2692 5804 2748
rect 5804 2692 5808 2748
rect 5744 2688 5808 2692
rect 5824 2748 5888 2752
rect 5824 2692 5828 2748
rect 5828 2692 5884 2748
rect 5884 2692 5888 2748
rect 5824 2688 5888 2692
rect 14848 2748 14912 2752
rect 14848 2692 14852 2748
rect 14852 2692 14908 2748
rect 14908 2692 14912 2748
rect 14848 2688 14912 2692
rect 14928 2748 14992 2752
rect 14928 2692 14932 2748
rect 14932 2692 14988 2748
rect 14988 2692 14992 2748
rect 14928 2688 14992 2692
rect 15008 2748 15072 2752
rect 15008 2692 15012 2748
rect 15012 2692 15068 2748
rect 15068 2692 15072 2748
rect 15008 2688 15072 2692
rect 15088 2748 15152 2752
rect 15088 2692 15092 2748
rect 15092 2692 15148 2748
rect 15148 2692 15152 2748
rect 15088 2688 15152 2692
rect 24112 2748 24176 2752
rect 24112 2692 24116 2748
rect 24116 2692 24172 2748
rect 24172 2692 24176 2748
rect 24112 2688 24176 2692
rect 24192 2748 24256 2752
rect 24192 2692 24196 2748
rect 24196 2692 24252 2748
rect 24252 2692 24256 2748
rect 24192 2688 24256 2692
rect 24272 2748 24336 2752
rect 24272 2692 24276 2748
rect 24276 2692 24332 2748
rect 24332 2692 24336 2748
rect 24272 2688 24336 2692
rect 24352 2748 24416 2752
rect 24352 2692 24356 2748
rect 24356 2692 24412 2748
rect 24412 2692 24416 2748
rect 24352 2688 24416 2692
rect 10216 2204 10280 2208
rect 10216 2148 10220 2204
rect 10220 2148 10276 2204
rect 10276 2148 10280 2204
rect 10216 2144 10280 2148
rect 10296 2204 10360 2208
rect 10296 2148 10300 2204
rect 10300 2148 10356 2204
rect 10356 2148 10360 2204
rect 10296 2144 10360 2148
rect 10376 2204 10440 2208
rect 10376 2148 10380 2204
rect 10380 2148 10436 2204
rect 10436 2148 10440 2204
rect 10376 2144 10440 2148
rect 10456 2204 10520 2208
rect 10456 2148 10460 2204
rect 10460 2148 10516 2204
rect 10516 2148 10520 2204
rect 10456 2144 10520 2148
rect 19480 2204 19544 2208
rect 19480 2148 19484 2204
rect 19484 2148 19540 2204
rect 19540 2148 19544 2204
rect 19480 2144 19544 2148
rect 19560 2204 19624 2208
rect 19560 2148 19564 2204
rect 19564 2148 19620 2204
rect 19620 2148 19624 2204
rect 19560 2144 19624 2148
rect 19640 2204 19704 2208
rect 19640 2148 19644 2204
rect 19644 2148 19700 2204
rect 19700 2148 19704 2204
rect 19640 2144 19704 2148
rect 19720 2204 19784 2208
rect 19720 2148 19724 2204
rect 19724 2148 19780 2204
rect 19780 2148 19784 2204
rect 19720 2144 19784 2148
<< metal4 >>
rect 5576 27776 5896 27792
rect 5576 27712 5584 27776
rect 5648 27712 5664 27776
rect 5728 27712 5744 27776
rect 5808 27712 5824 27776
rect 5888 27712 5896 27776
rect 5576 26688 5896 27712
rect 5576 26624 5584 26688
rect 5648 26624 5664 26688
rect 5728 26624 5744 26688
rect 5808 26624 5824 26688
rect 5888 26624 5896 26688
rect 5576 25600 5896 26624
rect 5576 25536 5584 25600
rect 5648 25536 5664 25600
rect 5728 25536 5744 25600
rect 5808 25536 5824 25600
rect 5888 25536 5896 25600
rect 5576 24512 5896 25536
rect 5576 24448 5584 24512
rect 5648 24448 5664 24512
rect 5728 24448 5744 24512
rect 5808 24448 5824 24512
rect 5888 24448 5896 24512
rect 5576 23424 5896 24448
rect 5576 23360 5584 23424
rect 5648 23360 5664 23424
rect 5728 23360 5744 23424
rect 5808 23360 5824 23424
rect 5888 23360 5896 23424
rect 5576 22336 5896 23360
rect 5576 22272 5584 22336
rect 5648 22272 5664 22336
rect 5728 22272 5744 22336
rect 5808 22272 5824 22336
rect 5888 22272 5896 22336
rect 5576 21248 5896 22272
rect 5576 21184 5584 21248
rect 5648 21184 5664 21248
rect 5728 21184 5744 21248
rect 5808 21184 5824 21248
rect 5888 21184 5896 21248
rect 5576 20160 5896 21184
rect 5576 20096 5584 20160
rect 5648 20096 5664 20160
rect 5728 20096 5744 20160
rect 5808 20096 5824 20160
rect 5888 20096 5896 20160
rect 5576 19072 5896 20096
rect 5576 19008 5584 19072
rect 5648 19008 5664 19072
rect 5728 19008 5744 19072
rect 5808 19008 5824 19072
rect 5888 19008 5896 19072
rect 5576 17984 5896 19008
rect 5576 17920 5584 17984
rect 5648 17920 5664 17984
rect 5728 17920 5744 17984
rect 5808 17920 5824 17984
rect 5888 17920 5896 17984
rect 5576 16896 5896 17920
rect 5576 16832 5584 16896
rect 5648 16832 5664 16896
rect 5728 16832 5744 16896
rect 5808 16832 5824 16896
rect 5888 16832 5896 16896
rect 5576 15808 5896 16832
rect 5576 15744 5584 15808
rect 5648 15744 5664 15808
rect 5728 15744 5744 15808
rect 5808 15744 5824 15808
rect 5888 15744 5896 15808
rect 5576 14720 5896 15744
rect 5576 14656 5584 14720
rect 5648 14656 5664 14720
rect 5728 14656 5744 14720
rect 5808 14656 5824 14720
rect 5888 14656 5896 14720
rect 5576 13632 5896 14656
rect 5576 13568 5584 13632
rect 5648 13568 5664 13632
rect 5728 13568 5744 13632
rect 5808 13568 5824 13632
rect 5888 13568 5896 13632
rect 5576 12544 5896 13568
rect 5576 12480 5584 12544
rect 5648 12480 5664 12544
rect 5728 12480 5744 12544
rect 5808 12480 5824 12544
rect 5888 12480 5896 12544
rect 5576 11456 5896 12480
rect 5576 11392 5584 11456
rect 5648 11392 5664 11456
rect 5728 11392 5744 11456
rect 5808 11392 5824 11456
rect 5888 11392 5896 11456
rect 5576 10368 5896 11392
rect 5576 10304 5584 10368
rect 5648 10304 5664 10368
rect 5728 10304 5744 10368
rect 5808 10304 5824 10368
rect 5888 10304 5896 10368
rect 5576 9280 5896 10304
rect 5576 9216 5584 9280
rect 5648 9216 5664 9280
rect 5728 9216 5744 9280
rect 5808 9216 5824 9280
rect 5888 9216 5896 9280
rect 5576 8192 5896 9216
rect 5576 8128 5584 8192
rect 5648 8128 5664 8192
rect 5728 8128 5744 8192
rect 5808 8128 5824 8192
rect 5888 8128 5896 8192
rect 5576 7104 5896 8128
rect 5576 7040 5584 7104
rect 5648 7040 5664 7104
rect 5728 7040 5744 7104
rect 5808 7040 5824 7104
rect 5888 7040 5896 7104
rect 5576 6016 5896 7040
rect 5576 5952 5584 6016
rect 5648 5952 5664 6016
rect 5728 5952 5744 6016
rect 5808 5952 5824 6016
rect 5888 5952 5896 6016
rect 5576 4928 5896 5952
rect 5576 4864 5584 4928
rect 5648 4864 5664 4928
rect 5728 4864 5744 4928
rect 5808 4864 5824 4928
rect 5888 4864 5896 4928
rect 5576 3840 5896 4864
rect 5576 3776 5584 3840
rect 5648 3776 5664 3840
rect 5728 3776 5744 3840
rect 5808 3776 5824 3840
rect 5888 3776 5896 3840
rect 5576 2752 5896 3776
rect 5576 2688 5584 2752
rect 5648 2688 5664 2752
rect 5728 2688 5744 2752
rect 5808 2688 5824 2752
rect 5888 2688 5896 2752
rect 5576 2128 5896 2688
rect 10208 27232 10528 27792
rect 10208 27168 10216 27232
rect 10280 27168 10296 27232
rect 10360 27168 10376 27232
rect 10440 27168 10456 27232
rect 10520 27168 10528 27232
rect 10208 26144 10528 27168
rect 10208 26080 10216 26144
rect 10280 26080 10296 26144
rect 10360 26080 10376 26144
rect 10440 26080 10456 26144
rect 10520 26080 10528 26144
rect 10208 25056 10528 26080
rect 10208 24992 10216 25056
rect 10280 24992 10296 25056
rect 10360 24992 10376 25056
rect 10440 24992 10456 25056
rect 10520 24992 10528 25056
rect 10208 23968 10528 24992
rect 10208 23904 10216 23968
rect 10280 23904 10296 23968
rect 10360 23904 10376 23968
rect 10440 23904 10456 23968
rect 10520 23904 10528 23968
rect 10208 22880 10528 23904
rect 10208 22816 10216 22880
rect 10280 22816 10296 22880
rect 10360 22816 10376 22880
rect 10440 22816 10456 22880
rect 10520 22816 10528 22880
rect 10208 21792 10528 22816
rect 10208 21728 10216 21792
rect 10280 21728 10296 21792
rect 10360 21728 10376 21792
rect 10440 21728 10456 21792
rect 10520 21728 10528 21792
rect 10208 20704 10528 21728
rect 10208 20640 10216 20704
rect 10280 20640 10296 20704
rect 10360 20640 10376 20704
rect 10440 20640 10456 20704
rect 10520 20640 10528 20704
rect 10208 19616 10528 20640
rect 10208 19552 10216 19616
rect 10280 19552 10296 19616
rect 10360 19552 10376 19616
rect 10440 19552 10456 19616
rect 10520 19552 10528 19616
rect 10208 18528 10528 19552
rect 10208 18464 10216 18528
rect 10280 18464 10296 18528
rect 10360 18464 10376 18528
rect 10440 18464 10456 18528
rect 10520 18464 10528 18528
rect 10208 17440 10528 18464
rect 10208 17376 10216 17440
rect 10280 17376 10296 17440
rect 10360 17376 10376 17440
rect 10440 17376 10456 17440
rect 10520 17376 10528 17440
rect 10208 16352 10528 17376
rect 14840 27776 15160 27792
rect 14840 27712 14848 27776
rect 14912 27712 14928 27776
rect 14992 27712 15008 27776
rect 15072 27712 15088 27776
rect 15152 27712 15160 27776
rect 14840 26688 15160 27712
rect 14840 26624 14848 26688
rect 14912 26624 14928 26688
rect 14992 26624 15008 26688
rect 15072 26624 15088 26688
rect 15152 26624 15160 26688
rect 14840 25600 15160 26624
rect 14840 25536 14848 25600
rect 14912 25536 14928 25600
rect 14992 25536 15008 25600
rect 15072 25536 15088 25600
rect 15152 25536 15160 25600
rect 14840 24512 15160 25536
rect 14840 24448 14848 24512
rect 14912 24448 14928 24512
rect 14992 24448 15008 24512
rect 15072 24448 15088 24512
rect 15152 24448 15160 24512
rect 14840 23424 15160 24448
rect 14840 23360 14848 23424
rect 14912 23360 14928 23424
rect 14992 23360 15008 23424
rect 15072 23360 15088 23424
rect 15152 23360 15160 23424
rect 14840 22336 15160 23360
rect 14840 22272 14848 22336
rect 14912 22272 14928 22336
rect 14992 22272 15008 22336
rect 15072 22272 15088 22336
rect 15152 22272 15160 22336
rect 14840 21248 15160 22272
rect 19472 27232 19792 27792
rect 19472 27168 19480 27232
rect 19544 27168 19560 27232
rect 19624 27168 19640 27232
rect 19704 27168 19720 27232
rect 19784 27168 19792 27232
rect 19472 26144 19792 27168
rect 19472 26080 19480 26144
rect 19544 26080 19560 26144
rect 19624 26080 19640 26144
rect 19704 26080 19720 26144
rect 19784 26080 19792 26144
rect 19472 25056 19792 26080
rect 19472 24992 19480 25056
rect 19544 24992 19560 25056
rect 19624 24992 19640 25056
rect 19704 24992 19720 25056
rect 19784 24992 19792 25056
rect 19472 23968 19792 24992
rect 19472 23904 19480 23968
rect 19544 23904 19560 23968
rect 19624 23904 19640 23968
rect 19704 23904 19720 23968
rect 19784 23904 19792 23968
rect 19472 22880 19792 23904
rect 19472 22816 19480 22880
rect 19544 22816 19560 22880
rect 19624 22816 19640 22880
rect 19704 22816 19720 22880
rect 19784 22816 19792 22880
rect 19472 21792 19792 22816
rect 19472 21728 19480 21792
rect 19544 21728 19560 21792
rect 19624 21728 19640 21792
rect 19704 21728 19720 21792
rect 19784 21728 19792 21792
rect 17539 21316 17605 21317
rect 17539 21252 17540 21316
rect 17604 21252 17605 21316
rect 17539 21251 17605 21252
rect 14840 21184 14848 21248
rect 14912 21184 14928 21248
rect 14992 21184 15008 21248
rect 15072 21184 15088 21248
rect 15152 21184 15160 21248
rect 14840 20160 15160 21184
rect 14840 20096 14848 20160
rect 14912 20096 14928 20160
rect 14992 20096 15008 20160
rect 15072 20096 15088 20160
rect 15152 20096 15160 20160
rect 14840 19072 15160 20096
rect 14840 19008 14848 19072
rect 14912 19008 14928 19072
rect 14992 19008 15008 19072
rect 15072 19008 15088 19072
rect 15152 19008 15160 19072
rect 14840 17984 15160 19008
rect 14840 17920 14848 17984
rect 14912 17920 14928 17984
rect 14992 17920 15008 17984
rect 15072 17920 15088 17984
rect 15152 17920 15160 17984
rect 14840 16896 15160 17920
rect 14840 16832 14848 16896
rect 14912 16832 14928 16896
rect 14992 16832 15008 16896
rect 15072 16832 15088 16896
rect 15152 16832 15160 16896
rect 13859 16692 13925 16693
rect 13859 16628 13860 16692
rect 13924 16628 13925 16692
rect 13859 16627 13925 16628
rect 14227 16692 14293 16693
rect 14227 16628 14228 16692
rect 14292 16628 14293 16692
rect 14227 16627 14293 16628
rect 10208 16288 10216 16352
rect 10280 16288 10296 16352
rect 10360 16288 10376 16352
rect 10440 16288 10456 16352
rect 10520 16288 10528 16352
rect 10208 15264 10528 16288
rect 10208 15200 10216 15264
rect 10280 15200 10296 15264
rect 10360 15200 10376 15264
rect 10440 15200 10456 15264
rect 10520 15200 10528 15264
rect 10208 14176 10528 15200
rect 10208 14112 10216 14176
rect 10280 14112 10296 14176
rect 10360 14112 10376 14176
rect 10440 14112 10456 14176
rect 10520 14112 10528 14176
rect 10208 13088 10528 14112
rect 10208 13024 10216 13088
rect 10280 13024 10296 13088
rect 10360 13024 10376 13088
rect 10440 13024 10456 13088
rect 10520 13024 10528 13088
rect 10208 12000 10528 13024
rect 10208 11936 10216 12000
rect 10280 11936 10296 12000
rect 10360 11936 10376 12000
rect 10440 11936 10456 12000
rect 10520 11936 10528 12000
rect 10208 10912 10528 11936
rect 11099 11116 11165 11117
rect 11099 11052 11100 11116
rect 11164 11052 11165 11116
rect 11099 11051 11165 11052
rect 10208 10848 10216 10912
rect 10280 10848 10296 10912
rect 10360 10848 10376 10912
rect 10440 10848 10456 10912
rect 10520 10848 10528 10912
rect 10208 9824 10528 10848
rect 10208 9760 10216 9824
rect 10280 9760 10296 9824
rect 10360 9760 10376 9824
rect 10440 9760 10456 9824
rect 10520 9760 10528 9824
rect 10208 8736 10528 9760
rect 10208 8672 10216 8736
rect 10280 8672 10296 8736
rect 10360 8672 10376 8736
rect 10440 8672 10456 8736
rect 10520 8672 10528 8736
rect 10208 7648 10528 8672
rect 11102 7989 11162 11051
rect 11099 7988 11165 7989
rect 11099 7924 11100 7988
rect 11164 7924 11165 7988
rect 11099 7923 11165 7924
rect 10208 7584 10216 7648
rect 10280 7584 10296 7648
rect 10360 7584 10376 7648
rect 10440 7584 10456 7648
rect 10520 7584 10528 7648
rect 10208 6560 10528 7584
rect 10208 6496 10216 6560
rect 10280 6496 10296 6560
rect 10360 6496 10376 6560
rect 10440 6496 10456 6560
rect 10520 6496 10528 6560
rect 10208 5472 10528 6496
rect 10208 5408 10216 5472
rect 10280 5408 10296 5472
rect 10360 5408 10376 5472
rect 10440 5408 10456 5472
rect 10520 5408 10528 5472
rect 10208 4384 10528 5408
rect 10208 4320 10216 4384
rect 10280 4320 10296 4384
rect 10360 4320 10376 4384
rect 10440 4320 10456 4384
rect 10520 4320 10528 4384
rect 10208 3296 10528 4320
rect 13862 3501 13922 16627
rect 14230 5949 14290 16627
rect 14840 15808 15160 16832
rect 14840 15744 14848 15808
rect 14912 15744 14928 15808
rect 14992 15744 15008 15808
rect 15072 15744 15088 15808
rect 15152 15744 15160 15808
rect 14840 14720 15160 15744
rect 14840 14656 14848 14720
rect 14912 14656 14928 14720
rect 14992 14656 15008 14720
rect 15072 14656 15088 14720
rect 15152 14656 15160 14720
rect 14840 13632 15160 14656
rect 15331 14516 15397 14517
rect 15331 14452 15332 14516
rect 15396 14452 15397 14516
rect 15331 14451 15397 14452
rect 14840 13568 14848 13632
rect 14912 13568 14928 13632
rect 14992 13568 15008 13632
rect 15072 13568 15088 13632
rect 15152 13568 15160 13632
rect 14840 12544 15160 13568
rect 15334 13293 15394 14451
rect 15331 13292 15397 13293
rect 15331 13228 15332 13292
rect 15396 13228 15397 13292
rect 15331 13227 15397 13228
rect 14840 12480 14848 12544
rect 14912 12480 14928 12544
rect 14992 12480 15008 12544
rect 15072 12480 15088 12544
rect 15152 12480 15160 12544
rect 14840 11456 15160 12480
rect 17542 12069 17602 21251
rect 19472 20704 19792 21728
rect 19472 20640 19480 20704
rect 19544 20640 19560 20704
rect 19624 20640 19640 20704
rect 19704 20640 19720 20704
rect 19784 20640 19792 20704
rect 19472 19616 19792 20640
rect 24104 27776 24424 27792
rect 24104 27712 24112 27776
rect 24176 27712 24192 27776
rect 24256 27712 24272 27776
rect 24336 27712 24352 27776
rect 24416 27712 24424 27776
rect 24104 26688 24424 27712
rect 24104 26624 24112 26688
rect 24176 26624 24192 26688
rect 24256 26624 24272 26688
rect 24336 26624 24352 26688
rect 24416 26624 24424 26688
rect 24104 25600 24424 26624
rect 24104 25536 24112 25600
rect 24176 25536 24192 25600
rect 24256 25536 24272 25600
rect 24336 25536 24352 25600
rect 24416 25536 24424 25600
rect 24104 24512 24424 25536
rect 24104 24448 24112 24512
rect 24176 24448 24192 24512
rect 24256 24448 24272 24512
rect 24336 24448 24352 24512
rect 24416 24448 24424 24512
rect 24104 23424 24424 24448
rect 24104 23360 24112 23424
rect 24176 23360 24192 23424
rect 24256 23360 24272 23424
rect 24336 23360 24352 23424
rect 24416 23360 24424 23424
rect 24104 22336 24424 23360
rect 24104 22272 24112 22336
rect 24176 22272 24192 22336
rect 24256 22272 24272 22336
rect 24336 22272 24352 22336
rect 24416 22272 24424 22336
rect 24104 21248 24424 22272
rect 24104 21184 24112 21248
rect 24176 21184 24192 21248
rect 24256 21184 24272 21248
rect 24336 21184 24352 21248
rect 24416 21184 24424 21248
rect 24104 20160 24424 21184
rect 24104 20096 24112 20160
rect 24176 20096 24192 20160
rect 24256 20096 24272 20160
rect 24336 20096 24352 20160
rect 24416 20096 24424 20160
rect 21035 19684 21101 19685
rect 21035 19620 21036 19684
rect 21100 19620 21101 19684
rect 21035 19619 21101 19620
rect 19472 19552 19480 19616
rect 19544 19552 19560 19616
rect 19624 19552 19640 19616
rect 19704 19552 19720 19616
rect 19784 19552 19792 19616
rect 19472 18528 19792 19552
rect 19472 18464 19480 18528
rect 19544 18464 19560 18528
rect 19624 18464 19640 18528
rect 19704 18464 19720 18528
rect 19784 18464 19792 18528
rect 19472 17440 19792 18464
rect 19472 17376 19480 17440
rect 19544 17376 19560 17440
rect 19624 17376 19640 17440
rect 19704 17376 19720 17440
rect 19784 17376 19792 17440
rect 19472 16352 19792 17376
rect 19472 16288 19480 16352
rect 19544 16288 19560 16352
rect 19624 16288 19640 16352
rect 19704 16288 19720 16352
rect 19784 16288 19792 16352
rect 19472 15264 19792 16288
rect 21038 15469 21098 19619
rect 24104 19072 24424 20096
rect 24104 19008 24112 19072
rect 24176 19008 24192 19072
rect 24256 19008 24272 19072
rect 24336 19008 24352 19072
rect 24416 19008 24424 19072
rect 24104 17984 24424 19008
rect 24104 17920 24112 17984
rect 24176 17920 24192 17984
rect 24256 17920 24272 17984
rect 24336 17920 24352 17984
rect 24416 17920 24424 17984
rect 24104 16896 24424 17920
rect 24104 16832 24112 16896
rect 24176 16832 24192 16896
rect 24256 16832 24272 16896
rect 24336 16832 24352 16896
rect 24416 16832 24424 16896
rect 24104 15808 24424 16832
rect 24104 15744 24112 15808
rect 24176 15744 24192 15808
rect 24256 15744 24272 15808
rect 24336 15744 24352 15808
rect 24416 15744 24424 15808
rect 21035 15468 21101 15469
rect 21035 15404 21036 15468
rect 21100 15404 21101 15468
rect 21035 15403 21101 15404
rect 19472 15200 19480 15264
rect 19544 15200 19560 15264
rect 19624 15200 19640 15264
rect 19704 15200 19720 15264
rect 19784 15200 19792 15264
rect 19472 14176 19792 15200
rect 19472 14112 19480 14176
rect 19544 14112 19560 14176
rect 19624 14112 19640 14176
rect 19704 14112 19720 14176
rect 19784 14112 19792 14176
rect 19472 13088 19792 14112
rect 19472 13024 19480 13088
rect 19544 13024 19560 13088
rect 19624 13024 19640 13088
rect 19704 13024 19720 13088
rect 19784 13024 19792 13088
rect 17539 12068 17605 12069
rect 17539 12004 17540 12068
rect 17604 12004 17605 12068
rect 17539 12003 17605 12004
rect 14840 11392 14848 11456
rect 14912 11392 14928 11456
rect 14992 11392 15008 11456
rect 15072 11392 15088 11456
rect 15152 11392 15160 11456
rect 14840 10368 15160 11392
rect 14840 10304 14848 10368
rect 14912 10304 14928 10368
rect 14992 10304 15008 10368
rect 15072 10304 15088 10368
rect 15152 10304 15160 10368
rect 14840 9280 15160 10304
rect 14840 9216 14848 9280
rect 14912 9216 14928 9280
rect 14992 9216 15008 9280
rect 15072 9216 15088 9280
rect 15152 9216 15160 9280
rect 14840 8192 15160 9216
rect 14840 8128 14848 8192
rect 14912 8128 14928 8192
rect 14992 8128 15008 8192
rect 15072 8128 15088 8192
rect 15152 8128 15160 8192
rect 14840 7104 15160 8128
rect 14840 7040 14848 7104
rect 14912 7040 14928 7104
rect 14992 7040 15008 7104
rect 15072 7040 15088 7104
rect 15152 7040 15160 7104
rect 14840 6016 15160 7040
rect 14840 5952 14848 6016
rect 14912 5952 14928 6016
rect 14992 5952 15008 6016
rect 15072 5952 15088 6016
rect 15152 5952 15160 6016
rect 14227 5948 14293 5949
rect 14227 5884 14228 5948
rect 14292 5884 14293 5948
rect 14227 5883 14293 5884
rect 14840 4928 15160 5952
rect 14840 4864 14848 4928
rect 14912 4864 14928 4928
rect 14992 4864 15008 4928
rect 15072 4864 15088 4928
rect 15152 4864 15160 4928
rect 14840 3840 15160 4864
rect 14840 3776 14848 3840
rect 14912 3776 14928 3840
rect 14992 3776 15008 3840
rect 15072 3776 15088 3840
rect 15152 3776 15160 3840
rect 13859 3500 13925 3501
rect 13859 3436 13860 3500
rect 13924 3436 13925 3500
rect 13859 3435 13925 3436
rect 10208 3232 10216 3296
rect 10280 3232 10296 3296
rect 10360 3232 10376 3296
rect 10440 3232 10456 3296
rect 10520 3232 10528 3296
rect 10208 2208 10528 3232
rect 10208 2144 10216 2208
rect 10280 2144 10296 2208
rect 10360 2144 10376 2208
rect 10440 2144 10456 2208
rect 10520 2144 10528 2208
rect 10208 2128 10528 2144
rect 14840 2752 15160 3776
rect 14840 2688 14848 2752
rect 14912 2688 14928 2752
rect 14992 2688 15008 2752
rect 15072 2688 15088 2752
rect 15152 2688 15160 2752
rect 14840 2128 15160 2688
rect 19472 12000 19792 13024
rect 19472 11936 19480 12000
rect 19544 11936 19560 12000
rect 19624 11936 19640 12000
rect 19704 11936 19720 12000
rect 19784 11936 19792 12000
rect 19472 10912 19792 11936
rect 19472 10848 19480 10912
rect 19544 10848 19560 10912
rect 19624 10848 19640 10912
rect 19704 10848 19720 10912
rect 19784 10848 19792 10912
rect 19472 9824 19792 10848
rect 19472 9760 19480 9824
rect 19544 9760 19560 9824
rect 19624 9760 19640 9824
rect 19704 9760 19720 9824
rect 19784 9760 19792 9824
rect 19472 8736 19792 9760
rect 19472 8672 19480 8736
rect 19544 8672 19560 8736
rect 19624 8672 19640 8736
rect 19704 8672 19720 8736
rect 19784 8672 19792 8736
rect 19472 7648 19792 8672
rect 19472 7584 19480 7648
rect 19544 7584 19560 7648
rect 19624 7584 19640 7648
rect 19704 7584 19720 7648
rect 19784 7584 19792 7648
rect 19472 6560 19792 7584
rect 19472 6496 19480 6560
rect 19544 6496 19560 6560
rect 19624 6496 19640 6560
rect 19704 6496 19720 6560
rect 19784 6496 19792 6560
rect 19472 5472 19792 6496
rect 19472 5408 19480 5472
rect 19544 5408 19560 5472
rect 19624 5408 19640 5472
rect 19704 5408 19720 5472
rect 19784 5408 19792 5472
rect 19472 4384 19792 5408
rect 19472 4320 19480 4384
rect 19544 4320 19560 4384
rect 19624 4320 19640 4384
rect 19704 4320 19720 4384
rect 19784 4320 19792 4384
rect 19472 3296 19792 4320
rect 19472 3232 19480 3296
rect 19544 3232 19560 3296
rect 19624 3232 19640 3296
rect 19704 3232 19720 3296
rect 19784 3232 19792 3296
rect 19472 2208 19792 3232
rect 19472 2144 19480 2208
rect 19544 2144 19560 2208
rect 19624 2144 19640 2208
rect 19704 2144 19720 2208
rect 19784 2144 19792 2208
rect 19472 2128 19792 2144
rect 24104 14720 24424 15744
rect 24104 14656 24112 14720
rect 24176 14656 24192 14720
rect 24256 14656 24272 14720
rect 24336 14656 24352 14720
rect 24416 14656 24424 14720
rect 24104 13632 24424 14656
rect 24104 13568 24112 13632
rect 24176 13568 24192 13632
rect 24256 13568 24272 13632
rect 24336 13568 24352 13632
rect 24416 13568 24424 13632
rect 24104 12544 24424 13568
rect 24104 12480 24112 12544
rect 24176 12480 24192 12544
rect 24256 12480 24272 12544
rect 24336 12480 24352 12544
rect 24416 12480 24424 12544
rect 24104 11456 24424 12480
rect 24104 11392 24112 11456
rect 24176 11392 24192 11456
rect 24256 11392 24272 11456
rect 24336 11392 24352 11456
rect 24416 11392 24424 11456
rect 24104 10368 24424 11392
rect 24104 10304 24112 10368
rect 24176 10304 24192 10368
rect 24256 10304 24272 10368
rect 24336 10304 24352 10368
rect 24416 10304 24424 10368
rect 24104 9280 24424 10304
rect 24104 9216 24112 9280
rect 24176 9216 24192 9280
rect 24256 9216 24272 9280
rect 24336 9216 24352 9280
rect 24416 9216 24424 9280
rect 24104 8192 24424 9216
rect 24104 8128 24112 8192
rect 24176 8128 24192 8192
rect 24256 8128 24272 8192
rect 24336 8128 24352 8192
rect 24416 8128 24424 8192
rect 24104 7104 24424 8128
rect 24104 7040 24112 7104
rect 24176 7040 24192 7104
rect 24256 7040 24272 7104
rect 24336 7040 24352 7104
rect 24416 7040 24424 7104
rect 24104 6016 24424 7040
rect 24104 5952 24112 6016
rect 24176 5952 24192 6016
rect 24256 5952 24272 6016
rect 24336 5952 24352 6016
rect 24416 5952 24424 6016
rect 24104 4928 24424 5952
rect 24104 4864 24112 4928
rect 24176 4864 24192 4928
rect 24256 4864 24272 4928
rect 24336 4864 24352 4928
rect 24416 4864 24424 4928
rect 24104 3840 24424 4864
rect 24104 3776 24112 3840
rect 24176 3776 24192 3840
rect 24256 3776 24272 3840
rect 24336 3776 24352 3840
rect 24416 3776 24424 3840
rect 24104 2752 24424 3776
rect 24104 2688 24112 2752
rect 24176 2688 24192 2752
rect 24256 2688 24272 2752
rect 24336 2688 24352 2752
rect 24416 2688 24424 2752
rect 24104 2128 24424 2688
use sky130_fd_sc_hd__diode_2  ANTENNA__0583__B pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 18216 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0583__C
timestamp 1644511149
transform 1 0 18676 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0584__A
timestamp 1644511149
transform 1 0 19228 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0585__A
timestamp 1644511149
transform 1 0 18952 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0585__B
timestamp 1644511149
transform 1 0 19872 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0585__C_N
timestamp 1644511149
transform 1 0 18308 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0586__A
timestamp 1644511149
transform -1 0 18676 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0587__B
timestamp 1644511149
transform 1 0 14628 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0593__B1
timestamp 1644511149
transform 1 0 16836 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0679__B1
timestamp 1644511149
transform 1 0 11500 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0693__A
timestamp 1644511149
transform -1 0 10580 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0696__A
timestamp 1644511149
transform -1 0 6992 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0699__A
timestamp 1644511149
transform 1 0 7636 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0702__A
timestamp 1644511149
transform 1 0 9752 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0722__C1
timestamp 1644511149
transform 1 0 11500 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0730__C1
timestamp 1644511149
transform 1 0 10948 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0734__A
timestamp 1644511149
transform 1 0 8188 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0740__C1
timestamp 1644511149
transform 1 0 9384 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0751__C1
timestamp 1644511149
transform 1 0 6532 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0756__B1
timestamp 1644511149
transform -1 0 8096 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0758__A_N
timestamp 1644511149
transform -1 0 19688 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0760__A
timestamp 1644511149
transform 1 0 18492 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0761__A
timestamp 1644511149
transform -1 0 24196 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0761__B
timestamp 1644511149
transform -1 0 24564 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0761__C
timestamp 1644511149
transform 1 0 23920 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0766__A
timestamp 1644511149
transform 1 0 16652 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0767__A
timestamp 1644511149
transform -1 0 18308 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0769__A_N
timestamp 1644511149
transform -1 0 15548 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0769__B
timestamp 1644511149
transform -1 0 18492 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0769__C
timestamp 1644511149
transform 1 0 15548 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0784__C1
timestamp 1644511149
transform 1 0 14996 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0791__C1
timestamp 1644511149
transform -1 0 14904 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0796__C1
timestamp 1644511149
transform -1 0 23000 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0801__C1
timestamp 1644511149
transform 1 0 16192 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0838__A0
timestamp 1644511149
transform 1 0 14168 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0842__A0
timestamp 1644511149
transform -1 0 17940 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0845__A0
timestamp 1644511149
transform 1 0 17112 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0848__A0
timestamp 1644511149
transform 1 0 17112 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0851__A0
timestamp 1644511149
transform 1 0 16008 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0854__A0
timestamp 1644511149
transform 1 0 14076 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0865__A
timestamp 1644511149
transform 1 0 18676 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0870__B1
timestamp 1644511149
transform 1 0 15824 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0879__B1
timestamp 1644511149
transform 1 0 17756 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0888__A
timestamp 1644511149
transform 1 0 17848 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0896__B1
timestamp 1644511149
transform 1 0 20240 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0900__A
timestamp 1644511149
transform 1 0 23184 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0911__A1
timestamp 1644511149
transform 1 0 13708 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0913__A1
timestamp 1644511149
transform 1 0 14904 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0915__A1
timestamp 1644511149
transform 1 0 17020 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0917__A1
timestamp 1644511149
transform 1 0 19228 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0919__A1
timestamp 1644511149
transform -1 0 14444 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0921__A1
timestamp 1644511149
transform 1 0 14536 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0924__A1
timestamp 1644511149
transform 1 0 13156 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0925__A_N
timestamp 1644511149
transform -1 0 13248 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0925__B
timestamp 1644511149
transform 1 0 12788 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0925__C
timestamp 1644511149
transform 1 0 17756 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0925__D
timestamp 1644511149
transform 1 0 16100 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0926__A
timestamp 1644511149
transform -1 0 15916 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0929__A
timestamp 1644511149
transform -1 0 21344 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0933__A0
timestamp 1644511149
transform 1 0 19688 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0936__A0
timestamp 1644511149
transform 1 0 20056 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0939__A0
timestamp 1644511149
transform 1 0 19228 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0942__A0
timestamp 1644511149
transform -1 0 21896 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0945__A0
timestamp 1644511149
transform 1 0 21344 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0949__A0
timestamp 1644511149
transform 1 0 15180 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0952__A0
timestamp 1644511149
transform 1 0 13156 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0955__A0
timestamp 1644511149
transform 1 0 16836 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0958__A
timestamp 1644511149
transform 1 0 12696 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0959__B
timestamp 1644511149
transform -1 0 24932 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0967__A1
timestamp 1644511149
transform -1 0 20608 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0969__A1
timestamp 1644511149
transform 1 0 21988 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0972__A1
timestamp 1644511149
transform 1 0 24380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0974__A1
timestamp 1644511149
transform 1 0 24656 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0976__A1
timestamp 1644511149
transform 1 0 25024 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0978__A1
timestamp 1644511149
transform -1 0 25300 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0980__A1
timestamp 1644511149
transform 1 0 25576 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1008__A
timestamp 1644511149
transform -1 0 24196 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1014__A0
timestamp 1644511149
transform 1 0 19320 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1017__A0
timestamp 1644511149
transform -1 0 25208 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1020__A0
timestamp 1644511149
transform -1 0 21160 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1023__A0
timestamp 1644511149
transform -1 0 26496 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1026__A0
timestamp 1644511149
transform -1 0 26220 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1029__A0
timestamp 1644511149
transform -1 0 21528 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1032__A0
timestamp 1644511149
transform -1 0 26588 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1046__B1
timestamp 1644511149
transform 1 0 20424 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1076__D
timestamp 1644511149
transform -1 0 8280 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1079__D
timestamp 1644511149
transform 1 0 8372 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clock_A
timestamp 1644511149
transform 1 0 12144 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_0_0_clock_A
timestamp 1644511149
transform -1 0 9660 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_1_0_clock_A
timestamp 1644511149
transform 1 0 12972 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_2_0_clock_A
timestamp 1644511149
transform 1 0 22172 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_3_0_clock_A
timestamp 1644511149
transform -1 0 24564 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_4_0_clock_A
timestamp 1644511149
transform 1 0 10580 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_5_0_clock_A
timestamp 1644511149
transform 1 0 10488 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_6_0_clock_A
timestamp 1644511149
transform 1 0 21068 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_7_0_clock_A
timestamp 1644511149
transform 1 0 19872 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1644511149
transform -1 0 1564 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1644511149
transform -1 0 2484 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1644511149
transform -1 0 11132 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1644511149
transform -1 0 27876 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1644511149
transform -1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1644511149
transform -1 0 27600 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1644511149
transform -1 0 1564 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1644511149
transform -1 0 27968 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1644511149
transform -1 0 21344 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1644511149
transform -1 0 2116 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1644511149
transform -1 0 27876 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1644511149
transform -1 0 1564 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1644511149
transform -1 0 5060 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1644511149
transform -1 0 27876 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1644511149
transform -1 0 16376 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1644511149
transform 1 0 23920 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1644511149
transform -1 0 22448 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1644511149
transform -1 0 2484 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1644511149
transform -1 0 2300 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1644511149
transform -1 0 2116 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1644511149
transform -1 0 27876 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9
timestamp 1644511149
transform 1 0 1932 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 4048 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40
timestamp 1644511149
transform 1 0 4784 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43
timestamp 1644511149
transform 1 0 5060 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 5796 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55
timestamp 1644511149
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57
timestamp 1644511149
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_62
timestamp 1644511149
transform 1 0 6808 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_74
timestamp 1644511149
transform 1 0 7912 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82
timestamp 1644511149
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_85
timestamp 1644511149
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_97
timestamp 1644511149
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_113
timestamp 1644511149
transform 1 0 11500 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_121
timestamp 1644511149
transform 1 0 12236 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_125
timestamp 1644511149
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1644511149
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_141
timestamp 1644511149
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_153
timestamp 1644511149
transform 1 0 15180 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_161
timestamp 1644511149
transform 1 0 15916 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_166
timestamp 1644511149
transform 1 0 16376 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169
timestamp 1644511149
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_177
timestamp 1644511149
transform 1 0 17388 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_189
timestamp 1644511149
transform 1 0 18492 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_194
timestamp 1644511149
transform 1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_207 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20148 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_216
timestamp 1644511149
transform 1 0 20976 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_220
timestamp 1644511149
transform 1 0 21344 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_225
timestamp 1644511149
transform 1 0 21804 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_231
timestamp 1644511149
transform 1 0 22356 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_243
timestamp 1644511149
transform 1 0 23460 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_251
timestamp 1644511149
transform 1 0 24196 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_253
timestamp 1644511149
transform 1 0 24380 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_261
timestamp 1644511149
transform 1 0 25116 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_266
timestamp 1644511149
transform 1 0 25576 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_278
timestamp 1644511149
transform 1 0 26680 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_284
timestamp 1644511149
transform 1 0 27232 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_288
timestamp 1644511149
transform 1 0 27600 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_294
timestamp 1644511149
transform 1 0 28152 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_298
timestamp 1644511149
transform 1 0 28520 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_5
timestamp 1644511149
transform 1 0 1564 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_17
timestamp 1644511149
transform 1 0 2668 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_29
timestamp 1644511149
transform 1 0 3772 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_41
timestamp 1644511149
transform 1 0 4876 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_53
timestamp 1644511149
transform 1 0 5980 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_57
timestamp 1644511149
transform 1 0 6348 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_74
timestamp 1644511149
transform 1 0 7912 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_78
timestamp 1644511149
transform 1 0 8280 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_90
timestamp 1644511149
transform 1 0 9384 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_102
timestamp 1644511149
transform 1 0 10488 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_110
timestamp 1644511149
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_113
timestamp 1644511149
transform 1 0 11500 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_131
timestamp 1644511149
transform 1 0 13156 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_149
timestamp 1644511149
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1644511149
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1644511149
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_169
timestamp 1644511149
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_181
timestamp 1644511149
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_193
timestamp 1644511149
transform 1 0 18860 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_210
timestamp 1644511149
transform 1 0 20424 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_222
timestamp 1644511149
transform 1 0 21528 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_225
timestamp 1644511149
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_237
timestamp 1644511149
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_249
timestamp 1644511149
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_261
timestamp 1644511149
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp 1644511149
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1644511149
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_281
timestamp 1644511149
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_297
timestamp 1644511149
transform 1 0 28428 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1644511149
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1644511149
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1644511149
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_29
timestamp 1644511149
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_41
timestamp 1644511149
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_53
timestamp 1644511149
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_65
timestamp 1644511149
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1644511149
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1644511149
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_85
timestamp 1644511149
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_97
timestamp 1644511149
transform 1 0 10028 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_105
timestamp 1644511149
transform 1 0 10764 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_110
timestamp 1644511149
transform 1 0 11224 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_117
timestamp 1644511149
transform 1 0 11868 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_123
timestamp 1644511149
transform 1 0 12420 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_127
timestamp 1644511149
transform 1 0 12788 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_132
timestamp 1644511149
transform 1 0 13248 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_138
timestamp 1644511149
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_141
timestamp 1644511149
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_153
timestamp 1644511149
transform 1 0 15180 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_161
timestamp 1644511149
transform 1 0 15916 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_180
timestamp 1644511149
transform 1 0 17664 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_188
timestamp 1644511149
transform 1 0 18400 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_203
timestamp 1644511149
transform 1 0 19780 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_210
timestamp 1644511149
transform 1 0 20424 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_229
timestamp 1644511149
transform 1 0 22172 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_241
timestamp 1644511149
transform 1 0 23276 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_249
timestamp 1644511149
transform 1 0 24012 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_269
timestamp 1644511149
transform 1 0 25852 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_281
timestamp 1644511149
transform 1 0 26956 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_293
timestamp 1644511149
transform 1 0 28060 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1644511149
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1644511149
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1644511149
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1644511149
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1644511149
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1644511149
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_57
timestamp 1644511149
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_69
timestamp 1644511149
transform 1 0 7452 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_77
timestamp 1644511149
transform 1 0 8188 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_95
timestamp 1644511149
transform 1 0 9844 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_104
timestamp 1644511149
transform 1 0 10672 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_113
timestamp 1644511149
transform 1 0 11500 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_117
timestamp 1644511149
transform 1 0 11868 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_126
timestamp 1644511149
transform 1 0 12696 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_3_137
timestamp 1644511149
transform 1 0 13708 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_156
timestamp 1644511149
transform 1 0 15456 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_173
timestamp 1644511149
transform 1 0 17020 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_178
timestamp 1644511149
transform 1 0 17480 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_190
timestamp 1644511149
transform 1 0 18584 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_200
timestamp 1644511149
transform 1 0 19504 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_3_222
timestamp 1644511149
transform 1 0 21528 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_232
timestamp 1644511149
transform 1 0 22448 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_252
timestamp 1644511149
transform 1 0 24288 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_264
timestamp 1644511149
transform 1 0 25392 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_276
timestamp 1644511149
transform 1 0 26496 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_281
timestamp 1644511149
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_293
timestamp 1644511149
transform 1 0 28060 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1644511149
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1644511149
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1644511149
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_29
timestamp 1644511149
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_41
timestamp 1644511149
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_53
timestamp 1644511149
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_65
timestamp 1644511149
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1644511149
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1644511149
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_85
timestamp 1644511149
transform 1 0 8924 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_4_96
timestamp 1644511149
transform 1 0 9936 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_115
timestamp 1644511149
transform 1 0 11684 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_127
timestamp 1644511149
transform 1 0 12788 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_135
timestamp 1644511149
transform 1 0 13524 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1644511149
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_151
timestamp 1644511149
transform 1 0 14996 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_158
timestamp 1644511149
transform 1 0 15640 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_162
timestamp 1644511149
transform 1 0 16008 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_170
timestamp 1644511149
transform 1 0 16744 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_178
timestamp 1644511149
transform 1 0 17480 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_186
timestamp 1644511149
transform 1 0 18216 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_193
timestamp 1644511149
transform 1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_204
timestamp 1644511149
transform 1 0 19872 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_210
timestamp 1644511149
transform 1 0 20424 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_218
timestamp 1644511149
transform 1 0 21160 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_226
timestamp 1644511149
transform 1 0 21896 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_232
timestamp 1644511149
transform 1 0 22448 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_239
timestamp 1644511149
transform 1 0 23092 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_244
timestamp 1644511149
transform 1 0 23552 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_253
timestamp 1644511149
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_265
timestamp 1644511149
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_277
timestamp 1644511149
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_289
timestamp 1644511149
transform 1 0 27692 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_293
timestamp 1644511149
transform 1 0 28060 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_297
timestamp 1644511149
transform 1 0 28428 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1644511149
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1644511149
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1644511149
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1644511149
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1644511149
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1644511149
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_57
timestamp 1644511149
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_69
timestamp 1644511149
transform 1 0 7452 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_73
timestamp 1644511149
transform 1 0 7820 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_90
timestamp 1644511149
transform 1 0 9384 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_96
timestamp 1644511149
transform 1 0 9936 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_102
timestamp 1644511149
transform 1 0 10488 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_108
timestamp 1644511149
transform 1 0 11040 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_120
timestamp 1644511149
transform 1 0 12144 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_127
timestamp 1644511149
transform 1 0 12788 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_134
timestamp 1644511149
transform 1 0 13432 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_140
timestamp 1644511149
transform 1 0 13984 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_146
timestamp 1644511149
transform 1 0 14536 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_155
timestamp 1644511149
transform 1 0 15364 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_166
timestamp 1644511149
transform 1 0 16376 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_185
timestamp 1644511149
transform 1 0 18124 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_197
timestamp 1644511149
transform 1 0 19228 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_204
timestamp 1644511149
transform 1 0 19872 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_216
timestamp 1644511149
transform 1 0 20976 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_225
timestamp 1644511149
transform 1 0 21804 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_231
timestamp 1644511149
transform 1 0 22356 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_237
timestamp 1644511149
transform 1 0 22908 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_242
timestamp 1644511149
transform 1 0 23368 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_262
timestamp 1644511149
transform 1 0 25208 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_274
timestamp 1644511149
transform 1 0 26312 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_5_281
timestamp 1644511149
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_293
timestamp 1644511149
transform 1 0 28060 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_6_7
timestamp 1644511149
transform 1 0 1748 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_19
timestamp 1644511149
transform 1 0 2852 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1644511149
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_29
timestamp 1644511149
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_41
timestamp 1644511149
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_53
timestamp 1644511149
transform 1 0 5980 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_77
timestamp 1644511149
transform 1 0 8188 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_81
timestamp 1644511149
transform 1 0 8556 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_85
timestamp 1644511149
transform 1 0 8924 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_90
timestamp 1644511149
transform 1 0 9384 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_99
timestamp 1644511149
transform 1 0 10212 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_103
timestamp 1644511149
transform 1 0 10580 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_111
timestamp 1644511149
transform 1 0 11316 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_121
timestamp 1644511149
transform 1 0 12236 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_127
timestamp 1644511149
transform 1 0 12788 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_131
timestamp 1644511149
transform 1 0 13156 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_138
timestamp 1644511149
transform 1 0 13800 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_141
timestamp 1644511149
transform 1 0 14076 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_151
timestamp 1644511149
transform 1 0 14996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_163
timestamp 1644511149
transform 1 0 16100 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_167
timestamp 1644511149
transform 1 0 16468 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_172
timestamp 1644511149
transform 1 0 16928 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_181
timestamp 1644511149
transform 1 0 17756 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_191
timestamp 1644511149
transform 1 0 18676 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1644511149
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_203
timestamp 1644511149
transform 1 0 19780 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_221
timestamp 1644511149
transform 1 0 21436 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_230
timestamp 1644511149
transform 1 0 22264 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_237
timestamp 1644511149
transform 1 0 22908 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_242
timestamp 1644511149
transform 1 0 23368 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_249
timestamp 1644511149
transform 1 0 24012 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_262
timestamp 1644511149
transform 1 0 25208 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_274
timestamp 1644511149
transform 1 0 26312 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_286
timestamp 1644511149
transform 1 0 27416 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_297
timestamp 1644511149
transform 1 0 28428 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1644511149
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1644511149
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1644511149
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1644511149
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1644511149
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1644511149
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_57
timestamp 1644511149
transform 1 0 6348 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_66
timestamp 1644511149
transform 1 0 7176 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_71
timestamp 1644511149
transform 1 0 7636 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_80
timestamp 1644511149
transform 1 0 8464 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_86
timestamp 1644511149
transform 1 0 9016 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_92
timestamp 1644511149
transform 1 0 9568 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_97
timestamp 1644511149
transform 1 0 10028 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_105
timestamp 1644511149
transform 1 0 10764 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_110
timestamp 1644511149
transform 1 0 11224 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_117
timestamp 1644511149
transform 1 0 11868 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_136
timestamp 1644511149
transform 1 0 13616 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_140
timestamp 1644511149
transform 1 0 13984 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_145
timestamp 1644511149
transform 1 0 14444 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_152
timestamp 1644511149
transform 1 0 15088 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_160
timestamp 1644511149
transform 1 0 15824 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_166
timestamp 1644511149
transform 1 0 16376 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_169
timestamp 1644511149
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_183
timestamp 1644511149
transform 1 0 17940 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_188
timestamp 1644511149
transform 1 0 18400 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_7_199
timestamp 1644511149
transform 1 0 19412 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_206
timestamp 1644511149
transform 1 0 20056 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_212
timestamp 1644511149
transform 1 0 20608 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_220
timestamp 1644511149
transform 1 0 21344 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_232
timestamp 1644511149
transform 1 0 22448 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_236
timestamp 1644511149
transform 1 0 22816 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_243
timestamp 1644511149
transform 1 0 23460 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_250
timestamp 1644511149
transform 1 0 24104 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_254
timestamp 1644511149
transform 1 0 24472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_259
timestamp 1644511149
transform 1 0 24932 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_268
timestamp 1644511149
transform 1 0 25760 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_281
timestamp 1644511149
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_293
timestamp 1644511149
transform 1 0 28060 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1644511149
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1644511149
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1644511149
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_29
timestamp 1644511149
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_41
timestamp 1644511149
transform 1 0 4876 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_61
timestamp 1644511149
transform 1 0 6716 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_68
timestamp 1644511149
transform 1 0 7360 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_79
timestamp 1644511149
transform 1 0 8372 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1644511149
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_101
timestamp 1644511149
transform 1 0 10396 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_110
timestamp 1644511149
transform 1 0 11224 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_115
timestamp 1644511149
transform 1 0 11684 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_124
timestamp 1644511149
transform 1 0 12512 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_130
timestamp 1644511149
transform 1 0 13064 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_138
timestamp 1644511149
transform 1 0 13800 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_157
timestamp 1644511149
transform 1 0 15548 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_175
timestamp 1644511149
transform 1 0 17204 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_181
timestamp 1644511149
transform 1 0 17756 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_192
timestamp 1644511149
transform 1 0 18768 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_200
timestamp 1644511149
transform 1 0 19504 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_208
timestamp 1644511149
transform 1 0 20240 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_212
timestamp 1644511149
transform 1 0 20608 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_221
timestamp 1644511149
transform 1 0 21436 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_227
timestamp 1644511149
transform 1 0 21988 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_231
timestamp 1644511149
transform 1 0 22356 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_250
timestamp 1644511149
transform 1 0 24104 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_253
timestamp 1644511149
transform 1 0 24380 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_260
timestamp 1644511149
transform 1 0 25024 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_278
timestamp 1644511149
transform 1 0 26680 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_290
timestamp 1644511149
transform 1 0 27784 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_298
timestamp 1644511149
transform 1 0 28520 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1644511149
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1644511149
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_27
timestamp 1644511149
transform 1 0 3588 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_35
timestamp 1644511149
transform 1 0 4324 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_54
timestamp 1644511149
transform 1 0 6072 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_67
timestamp 1644511149
transform 1 0 7268 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_76
timestamp 1644511149
transform 1 0 8096 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_80
timestamp 1644511149
transform 1 0 8464 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_85
timestamp 1644511149
transform 1 0 8924 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_91
timestamp 1644511149
transform 1 0 9476 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_97
timestamp 1644511149
transform 1 0 10028 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_110
timestamp 1644511149
transform 1 0 11224 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_113
timestamp 1644511149
transform 1 0 11500 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_119
timestamp 1644511149
transform 1 0 12052 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_131
timestamp 1644511149
transform 1 0 13156 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_143
timestamp 1644511149
transform 1 0 14260 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_9_153
timestamp 1644511149
transform 1 0 15180 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_159
timestamp 1644511149
transform 1 0 15732 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_164
timestamp 1644511149
transform 1 0 16192 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_169
timestamp 1644511149
transform 1 0 16652 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_9_179
timestamp 1644511149
transform 1 0 17572 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_197
timestamp 1644511149
transform 1 0 19228 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_211
timestamp 1644511149
transform 1 0 20516 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1644511149
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1644511149
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_231
timestamp 1644511149
transform 1 0 22356 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_239
timestamp 1644511149
transform 1 0 23092 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_245
timestamp 1644511149
transform 1 0 23644 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_249
timestamp 1644511149
transform 1 0 24012 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_259
timestamp 1644511149
transform 1 0 24932 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_266
timestamp 1644511149
transform 1 0 25576 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_278
timestamp 1644511149
transform 1 0 26680 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_281
timestamp 1644511149
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_293
timestamp 1644511149
transform 1 0 28060 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_10_5
timestamp 1644511149
transform 1 0 1564 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_17
timestamp 1644511149
transform 1 0 2668 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_25
timestamp 1644511149
transform 1 0 3404 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_29
timestamp 1644511149
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_41
timestamp 1644511149
transform 1 0 4876 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_49
timestamp 1644511149
transform 1 0 5612 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_55
timestamp 1644511149
transform 1 0 6164 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_65
timestamp 1644511149
transform 1 0 7084 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_69
timestamp 1644511149
transform 1 0 7452 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_73
timestamp 1644511149
transform 1 0 7820 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_78
timestamp 1644511149
transform 1 0 8280 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_10_85
timestamp 1644511149
transform 1 0 8924 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_10_93
timestamp 1644511149
transform 1 0 9660 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_99
timestamp 1644511149
transform 1 0 10212 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_108
timestamp 1644511149
transform 1 0 11040 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_112
timestamp 1644511149
transform 1 0 11408 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_119
timestamp 1644511149
transform 1 0 12052 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_125
timestamp 1644511149
transform 1 0 12604 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_135
timestamp 1644511149
transform 1 0 13524 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1644511149
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_146
timestamp 1644511149
transform 1 0 14536 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_10_158
timestamp 1644511149
transform 1 0 15640 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_162
timestamp 1644511149
transform 1 0 16008 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_169
timestamp 1644511149
transform 1 0 16652 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_178
timestamp 1644511149
transform 1 0 17480 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_184
timestamp 1644511149
transform 1 0 18032 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_188
timestamp 1644511149
transform 1 0 18400 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_194
timestamp 1644511149
transform 1 0 18952 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_204
timestamp 1644511149
transform 1 0 19872 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_212
timestamp 1644511149
transform 1 0 20608 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_221
timestamp 1644511149
transform 1 0 21436 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_239
timestamp 1644511149
transform 1 0 23092 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_243
timestamp 1644511149
transform 1 0 23460 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_247
timestamp 1644511149
transform 1 0 23828 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1644511149
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_256
timestamp 1644511149
transform 1 0 24656 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_262
timestamp 1644511149
transform 1 0 25208 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_272
timestamp 1644511149
transform 1 0 26128 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_284
timestamp 1644511149
transform 1 0 27232 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_10_292
timestamp 1644511149
transform 1 0 27968 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_297
timestamp 1644511149
transform 1 0 28428 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_3
timestamp 1644511149
transform 1 0 1380 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_11
timestamp 1644511149
transform 1 0 2116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_23
timestamp 1644511149
transform 1 0 3220 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_35
timestamp 1644511149
transform 1 0 4324 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_54
timestamp 1644511149
transform 1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_57
timestamp 1644511149
transform 1 0 6348 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_61
timestamp 1644511149
transform 1 0 6716 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_66
timestamp 1644511149
transform 1 0 7176 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_70
timestamp 1644511149
transform 1 0 7544 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_77
timestamp 1644511149
transform 1 0 8188 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_95
timestamp 1644511149
transform 1 0 9844 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_103
timestamp 1644511149
transform 1 0 10580 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_110
timestamp 1644511149
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_117
timestamp 1644511149
transform 1 0 11868 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_123
timestamp 1644511149
transform 1 0 12420 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_11_135
timestamp 1644511149
transform 1 0 13524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_11_148
timestamp 1644511149
transform 1 0 14720 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_166
timestamp 1644511149
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_174
timestamp 1644511149
transform 1 0 17112 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_181
timestamp 1644511149
transform 1 0 17756 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_186
timestamp 1644511149
transform 1 0 18216 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_190
timestamp 1644511149
transform 1 0 18584 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_193
timestamp 1644511149
transform 1 0 18860 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_199
timestamp 1644511149
transform 1 0 19412 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_11_218
timestamp 1644511149
transform 1 0 21160 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_11_225
timestamp 1644511149
transform 1 0 21804 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_231
timestamp 1644511149
transform 1 0 22356 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_237
timestamp 1644511149
transform 1 0 22908 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_11_259
timestamp 1644511149
transform 1 0 24932 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_278
timestamp 1644511149
transform 1 0 26680 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_281
timestamp 1644511149
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_293
timestamp 1644511149
transform 1 0 28060 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1644511149
transform 1 0 1380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_9
timestamp 1644511149
transform 1 0 1932 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_13
timestamp 1644511149
transform 1 0 2300 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_25
timestamp 1644511149
transform 1 0 3404 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_29
timestamp 1644511149
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_41
timestamp 1644511149
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_69
timestamp 1644511149
transform 1 0 7452 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1644511149
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1644511149
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_85
timestamp 1644511149
transform 1 0 8924 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_93
timestamp 1644511149
transform 1 0 9660 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_100
timestamp 1644511149
transform 1 0 10304 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_12_111
timestamp 1644511149
transform 1 0 11316 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_118
timestamp 1644511149
transform 1 0 11960 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_136
timestamp 1644511149
transform 1 0 13616 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_141
timestamp 1644511149
transform 1 0 14076 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_149
timestamp 1644511149
transform 1 0 14812 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_155
timestamp 1644511149
transform 1 0 15364 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_167
timestamp 1644511149
transform 1 0 16468 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_176
timestamp 1644511149
transform 1 0 17296 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_194
timestamp 1644511149
transform 1 0 18952 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_197
timestamp 1644511149
transform 1 0 19228 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_200
timestamp 1644511149
transform 1 0 19504 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_207
timestamp 1644511149
transform 1 0 20148 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_212
timestamp 1644511149
transform 1 0 20608 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_220
timestamp 1644511149
transform 1 0 21344 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_229
timestamp 1644511149
transform 1 0 22172 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_241
timestamp 1644511149
transform 1 0 23276 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_249
timestamp 1644511149
transform 1 0 24012 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_253
timestamp 1644511149
transform 1 0 24380 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_257
timestamp 1644511149
transform 1 0 24748 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_267
timestamp 1644511149
transform 1 0 25668 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_272
timestamp 1644511149
transform 1 0 26128 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_284
timestamp 1644511149
transform 1 0 27232 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_292
timestamp 1644511149
transform 1 0 27968 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_297
timestamp 1644511149
transform 1 0 28428 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1644511149
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1644511149
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1644511149
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_39
timestamp 1644511149
transform 1 0 4692 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_45
timestamp 1644511149
transform 1 0 5244 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_52
timestamp 1644511149
transform 1 0 5888 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_57
timestamp 1644511149
transform 1 0 6348 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_63
timestamp 1644511149
transform 1 0 6900 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_70
timestamp 1644511149
transform 1 0 7544 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_76
timestamp 1644511149
transform 1 0 8096 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_83
timestamp 1644511149
transform 1 0 8740 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_89
timestamp 1644511149
transform 1 0 9292 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_107
timestamp 1644511149
transform 1 0 10948 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1644511149
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_113
timestamp 1644511149
transform 1 0 11500 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_122
timestamp 1644511149
transform 1 0 12328 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_128
timestamp 1644511149
transform 1 0 12880 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_143
timestamp 1644511149
transform 1 0 14260 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_149
timestamp 1644511149
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_161
timestamp 1644511149
transform 1 0 15916 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_166
timestamp 1644511149
transform 1 0 16376 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_172
timestamp 1644511149
transform 1 0 16928 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_180
timestamp 1644511149
transform 1 0 17664 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_200
timestamp 1644511149
transform 1 0 19504 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_213
timestamp 1644511149
transform 1 0 20700 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_217
timestamp 1644511149
transform 1 0 21068 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_222
timestamp 1644511149
transform 1 0 21528 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_241
timestamp 1644511149
transform 1 0 23276 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_254
timestamp 1644511149
transform 1 0 24472 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_265
timestamp 1644511149
transform 1 0 25484 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_276
timestamp 1644511149
transform 1 0 26496 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_281
timestamp 1644511149
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_293
timestamp 1644511149
transform 1 0 28060 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1644511149
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1644511149
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1644511149
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_29
timestamp 1644511149
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_41
timestamp 1644511149
transform 1 0 4876 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_60
timestamp 1644511149
transform 1 0 6624 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_68
timestamp 1644511149
transform 1 0 7360 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_80
timestamp 1644511149
transform 1 0 8464 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_92
timestamp 1644511149
transform 1 0 9568 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_104
timestamp 1644511149
transform 1 0 10672 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_108
timestamp 1644511149
transform 1 0 11040 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_119
timestamp 1644511149
transform 1 0 12052 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_125
timestamp 1644511149
transform 1 0 12604 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_132
timestamp 1644511149
transform 1 0 13248 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_137
timestamp 1644511149
transform 1 0 13708 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_144
timestamp 1644511149
transform 1 0 14352 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_151
timestamp 1644511149
transform 1 0 14996 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_160
timestamp 1644511149
transform 1 0 15824 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_175
timestamp 1644511149
transform 1 0 17204 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_183
timestamp 1644511149
transform 1 0 17940 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_189
timestamp 1644511149
transform 1 0 18492 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_193
timestamp 1644511149
transform 1 0 18860 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_197
timestamp 1644511149
transform 1 0 19228 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_201
timestamp 1644511149
transform 1 0 19596 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_219
timestamp 1644511149
transform 1 0 21252 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_232
timestamp 1644511149
transform 1 0 22448 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_250
timestamp 1644511149
transform 1 0 24104 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_262
timestamp 1644511149
transform 1 0 25208 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_282
timestamp 1644511149
transform 1 0 27048 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_287
timestamp 1644511149
transform 1 0 27508 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_6
timestamp 1644511149
transform 1 0 1656 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_18
timestamp 1644511149
transform 1 0 2760 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_30
timestamp 1644511149
transform 1 0 3864 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_42
timestamp 1644511149
transform 1 0 4968 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_46
timestamp 1644511149
transform 1 0 5336 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_50
timestamp 1644511149
transform 1 0 5704 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_15_57
timestamp 1644511149
transform 1 0 6348 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_63
timestamp 1644511149
transform 1 0 6900 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_70
timestamp 1644511149
transform 1 0 7544 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_75
timestamp 1644511149
transform 1 0 8004 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_79
timestamp 1644511149
transform 1 0 8372 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_85
timestamp 1644511149
transform 1 0 8924 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_103
timestamp 1644511149
transform 1 0 10580 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_108
timestamp 1644511149
transform 1 0 11040 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_129
timestamp 1644511149
transform 1 0 12972 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_141
timestamp 1644511149
transform 1 0 14076 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_148
timestamp 1644511149
transform 1 0 14720 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_158
timestamp 1644511149
transform 1 0 15640 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_166
timestamp 1644511149
transform 1 0 16376 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_169
timestamp 1644511149
transform 1 0 16652 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_175
timestamp 1644511149
transform 1 0 17204 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_194
timestamp 1644511149
transform 1 0 18952 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_200
timestamp 1644511149
transform 1 0 19504 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_207
timestamp 1644511149
transform 1 0 20148 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_214
timestamp 1644511149
transform 1 0 20792 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_218
timestamp 1644511149
transform 1 0 21160 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_222
timestamp 1644511149
transform 1 0 21528 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_225
timestamp 1644511149
transform 1 0 21804 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_236
timestamp 1644511149
transform 1 0 22816 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_241
timestamp 1644511149
transform 1 0 23276 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_259
timestamp 1644511149
transform 1 0 24932 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_263
timestamp 1644511149
transform 1 0 25300 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_273
timestamp 1644511149
transform 1 0 26220 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_278
timestamp 1644511149
transform 1 0 26680 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_281
timestamp 1644511149
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_297
timestamp 1644511149
transform 1 0 28428 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1644511149
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1644511149
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1644511149
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_29
timestamp 1644511149
transform 1 0 3772 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_16_53
timestamp 1644511149
transform 1 0 5980 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_61
timestamp 1644511149
transform 1 0 6716 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_68
timestamp 1644511149
transform 1 0 7360 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_73
timestamp 1644511149
transform 1 0 7820 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_82
timestamp 1644511149
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_89
timestamp 1644511149
transform 1 0 9292 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_97
timestamp 1644511149
transform 1 0 10028 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_16_111
timestamp 1644511149
transform 1 0 11316 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_117
timestamp 1644511149
transform 1 0 11868 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_128
timestamp 1644511149
transform 1 0 12880 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_137
timestamp 1644511149
transform 1 0 13708 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_145
timestamp 1644511149
transform 1 0 14444 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_154
timestamp 1644511149
transform 1 0 15272 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_158
timestamp 1644511149
transform 1 0 15640 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_161
timestamp 1644511149
transform 1 0 15916 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_165
timestamp 1644511149
transform 1 0 16284 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_171
timestamp 1644511149
transform 1 0 16836 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_175
timestamp 1644511149
transform 1 0 17204 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_193
timestamp 1644511149
transform 1 0 18860 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_199
timestamp 1644511149
transform 1 0 19412 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_217
timestamp 1644511149
transform 1 0 21068 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_236
timestamp 1644511149
transform 1 0 22816 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_248
timestamp 1644511149
transform 1 0 23920 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_255
timestamp 1644511149
transform 1 0 24564 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_266
timestamp 1644511149
transform 1 0 25576 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_284
timestamp 1644511149
transform 1 0 27232 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_296
timestamp 1644511149
transform 1 0 28336 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1644511149
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1644511149
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_27
timestamp 1644511149
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_39
timestamp 1644511149
transform 1 0 4692 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_43
timestamp 1644511149
transform 1 0 5060 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_47
timestamp 1644511149
transform 1 0 5428 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_53
timestamp 1644511149
transform 1 0 5980 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_57
timestamp 1644511149
transform 1 0 6348 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_67
timestamp 1644511149
transform 1 0 7268 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_71
timestamp 1644511149
transform 1 0 7636 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_82
timestamp 1644511149
transform 1 0 8648 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_92
timestamp 1644511149
transform 1 0 9568 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_97
timestamp 1644511149
transform 1 0 10028 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_107
timestamp 1644511149
transform 1 0 10948 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1644511149
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_115
timestamp 1644511149
transform 1 0 11684 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_122
timestamp 1644511149
transform 1 0 12328 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_127
timestamp 1644511149
transform 1 0 12788 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_131
timestamp 1644511149
transform 1 0 13156 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_17_139
timestamp 1644511149
transform 1 0 13892 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_157
timestamp 1644511149
transform 1 0 15548 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_163
timestamp 1644511149
transform 1 0 16100 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1644511149
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_185
timestamp 1644511149
transform 1 0 18124 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_189
timestamp 1644511149
transform 1 0 18492 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_195
timestamp 1644511149
transform 1 0 19044 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_201
timestamp 1644511149
transform 1 0 19596 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_205
timestamp 1644511149
transform 1 0 19964 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_215
timestamp 1644511149
transform 1 0 20884 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_220
timestamp 1644511149
transform 1 0 21344 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_225
timestamp 1644511149
transform 1 0 21804 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_231
timestamp 1644511149
transform 1 0 22356 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_236
timestamp 1644511149
transform 1 0 22816 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_241
timestamp 1644511149
transform 1 0 23276 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_247
timestamp 1644511149
transform 1 0 23828 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_17_259
timestamp 1644511149
transform 1 0 24932 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_265
timestamp 1644511149
transform 1 0 25484 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_275
timestamp 1644511149
transform 1 0 26404 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1644511149
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_281
timestamp 1644511149
transform 1 0 26956 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_291
timestamp 1644511149
transform 1 0 27876 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_297
timestamp 1644511149
transform 1 0 28428 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1644511149
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1644511149
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1644511149
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_29
timestamp 1644511149
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_41
timestamp 1644511149
transform 1 0 4876 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_47
timestamp 1644511149
transform 1 0 5428 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_56
timestamp 1644511149
transform 1 0 6256 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_64
timestamp 1644511149
transform 1 0 6992 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_72
timestamp 1644511149
transform 1 0 7728 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_76
timestamp 1644511149
transform 1 0 8096 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_82
timestamp 1644511149
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_90
timestamp 1644511149
transform 1 0 9384 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_18_101
timestamp 1644511149
transform 1 0 10396 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_119
timestamp 1644511149
transform 1 0 12052 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_138
timestamp 1644511149
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_141
timestamp 1644511149
transform 1 0 14076 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_150
timestamp 1644511149
transform 1 0 14904 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_160
timestamp 1644511149
transform 1 0 15824 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_169
timestamp 1644511149
transform 1 0 16652 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_173
timestamp 1644511149
transform 1 0 17020 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_182
timestamp 1644511149
transform 1 0 17848 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_187
timestamp 1644511149
transform 1 0 18308 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_191
timestamp 1644511149
transform 1 0 18676 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1644511149
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_199
timestamp 1644511149
transform 1 0 19412 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_205
timestamp 1644511149
transform 1 0 19964 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_209
timestamp 1644511149
transform 1 0 20332 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_219
timestamp 1644511149
transform 1 0 21252 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_227
timestamp 1644511149
transform 1 0 21988 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_238
timestamp 1644511149
transform 1 0 23000 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_245
timestamp 1644511149
transform 1 0 23644 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_250
timestamp 1644511149
transform 1 0 24104 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_258
timestamp 1644511149
transform 1 0 24840 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_262
timestamp 1644511149
transform 1 0 25208 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_280
timestamp 1644511149
transform 1 0 26864 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_292
timestamp 1644511149
transform 1 0 27968 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_298
timestamp 1644511149
transform 1 0 28520 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1644511149
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1644511149
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_27
timestamp 1644511149
transform 1 0 3588 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_35
timestamp 1644511149
transform 1 0 4324 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_52
timestamp 1644511149
transform 1 0 5888 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_57
timestamp 1644511149
transform 1 0 6348 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_61
timestamp 1644511149
transform 1 0 6716 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_67
timestamp 1644511149
transform 1 0 7268 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_72
timestamp 1644511149
transform 1 0 7728 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_81
timestamp 1644511149
transform 1 0 8556 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_88
timestamp 1644511149
transform 1 0 9200 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_92
timestamp 1644511149
transform 1 0 9568 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_103
timestamp 1644511149
transform 1 0 10580 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_19_109
timestamp 1644511149
transform 1 0 11132 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_19_120
timestamp 1644511149
transform 1 0 12144 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_128
timestamp 1644511149
transform 1 0 12880 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_133
timestamp 1644511149
transform 1 0 13340 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_140
timestamp 1644511149
transform 1 0 13984 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_147
timestamp 1644511149
transform 1 0 14628 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_154
timestamp 1644511149
transform 1 0 15272 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_159
timestamp 1644511149
transform 1 0 15732 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_166
timestamp 1644511149
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_169
timestamp 1644511149
transform 1 0 16652 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_175
timestamp 1644511149
transform 1 0 17204 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_182
timestamp 1644511149
transform 1 0 17848 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_189
timestamp 1644511149
transform 1 0 18492 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_197
timestamp 1644511149
transform 1 0 19228 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_204
timestamp 1644511149
transform 1 0 19872 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_222
timestamp 1644511149
transform 1 0 21528 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_229
timestamp 1644511149
transform 1 0 22172 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_247
timestamp 1644511149
transform 1 0 23828 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_251
timestamp 1644511149
transform 1 0 24196 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_262
timestamp 1644511149
transform 1 0 25208 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_267
timestamp 1644511149
transform 1 0 25668 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_272
timestamp 1644511149
transform 1 0 26128 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_276
timestamp 1644511149
transform 1 0 26496 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_281
timestamp 1644511149
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_293
timestamp 1644511149
transform 1 0 28060 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_297
timestamp 1644511149
transform 1 0 28428 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1644511149
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1644511149
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1644511149
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_29
timestamp 1644511149
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_41
timestamp 1644511149
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_53
timestamp 1644511149
transform 1 0 5980 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_64
timestamp 1644511149
transform 1 0 6992 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_71
timestamp 1644511149
transform 1 0 7636 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_82
timestamp 1644511149
transform 1 0 8648 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_93
timestamp 1644511149
transform 1 0 9660 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_100
timestamp 1644511149
transform 1 0 10304 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_104
timestamp 1644511149
transform 1 0 10672 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_112
timestamp 1644511149
transform 1 0 11408 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_120
timestamp 1644511149
transform 1 0 12144 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_131
timestamp 1644511149
transform 1 0 13156 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_136
timestamp 1644511149
transform 1 0 13616 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_144
timestamp 1644511149
transform 1 0 14352 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_148
timestamp 1644511149
transform 1 0 14720 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_152
timestamp 1644511149
transform 1 0 15088 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_157
timestamp 1644511149
transform 1 0 15548 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_162
timestamp 1644511149
transform 1 0 16008 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_170
timestamp 1644511149
transform 1 0 16744 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_174
timestamp 1644511149
transform 1 0 17112 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_183
timestamp 1644511149
transform 1 0 17940 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_194
timestamp 1644511149
transform 1 0 18952 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_207
timestamp 1644511149
transform 1 0 20148 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_214
timestamp 1644511149
transform 1 0 20792 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_220
timestamp 1644511149
transform 1 0 21344 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_225
timestamp 1644511149
transform 1 0 21804 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_238
timestamp 1644511149
transform 1 0 23000 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_242
timestamp 1644511149
transform 1 0 23368 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_248
timestamp 1644511149
transform 1 0 23920 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_253
timestamp 1644511149
transform 1 0 24380 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_263
timestamp 1644511149
transform 1 0 25300 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_281
timestamp 1644511149
transform 1 0 26956 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_293
timestamp 1644511149
transform 1 0 28060 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_21_6
timestamp 1644511149
transform 1 0 1656 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_18
timestamp 1644511149
transform 1 0 2760 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_30
timestamp 1644511149
transform 1 0 3864 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_54
timestamp 1644511149
transform 1 0 6072 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_57
timestamp 1644511149
transform 1 0 6348 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_61
timestamp 1644511149
transform 1 0 6716 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_66
timestamp 1644511149
transform 1 0 7176 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_71
timestamp 1644511149
transform 1 0 7636 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_83
timestamp 1644511149
transform 1 0 8740 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_89
timestamp 1644511149
transform 1 0 9292 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_107
timestamp 1644511149
transform 1 0 10948 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1644511149
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_113
timestamp 1644511149
transform 1 0 11500 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_118
timestamp 1644511149
transform 1 0 11960 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_128
timestamp 1644511149
transform 1 0 12880 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_132
timestamp 1644511149
transform 1 0 13248 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_142
timestamp 1644511149
transform 1 0 14168 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_160
timestamp 1644511149
transform 1 0 15824 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_166
timestamp 1644511149
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_179
timestamp 1644511149
transform 1 0 17572 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_186
timestamp 1644511149
transform 1 0 18216 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_191
timestamp 1644511149
transform 1 0 18676 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_197
timestamp 1644511149
transform 1 0 19228 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_202
timestamp 1644511149
transform 1 0 19688 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_208
timestamp 1644511149
transform 1 0 20240 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_213
timestamp 1644511149
transform 1 0 20700 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_219
timestamp 1644511149
transform 1 0 21252 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1644511149
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_241
timestamp 1644511149
transform 1 0 23276 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_21_254
timestamp 1644511149
transform 1 0 24472 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_262
timestamp 1644511149
transform 1 0 25208 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_269
timestamp 1644511149
transform 1 0 25852 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_273
timestamp 1644511149
transform 1 0 26220 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_277
timestamp 1644511149
transform 1 0 26588 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_281
timestamp 1644511149
transform 1 0 26956 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_291
timestamp 1644511149
transform 1 0 27876 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_297
timestamp 1644511149
transform 1 0 28428 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1644511149
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1644511149
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1644511149
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_29
timestamp 1644511149
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_41
timestamp 1644511149
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_53
timestamp 1644511149
transform 1 0 5980 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_22_75
timestamp 1644511149
transform 1 0 8004 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1644511149
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_88
timestamp 1644511149
transform 1 0 9200 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_92
timestamp 1644511149
transform 1 0 9568 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_104
timestamp 1644511149
transform 1 0 10672 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_110
timestamp 1644511149
transform 1 0 11224 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_127
timestamp 1644511149
transform 1 0 12788 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_133
timestamp 1644511149
transform 1 0 13340 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_138
timestamp 1644511149
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_149
timestamp 1644511149
transform 1 0 14812 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_157
timestamp 1644511149
transform 1 0 15548 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_22_166
timestamp 1644511149
transform 1 0 16376 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_178
timestamp 1644511149
transform 1 0 17480 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_188
timestamp 1644511149
transform 1 0 18400 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_193
timestamp 1644511149
transform 1 0 18860 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_203
timestamp 1644511149
transform 1 0 19780 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_210
timestamp 1644511149
transform 1 0 20424 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_216
timestamp 1644511149
transform 1 0 20976 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_222
timestamp 1644511149
transform 1 0 21528 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_230
timestamp 1644511149
transform 1 0 22264 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_235
timestamp 1644511149
transform 1 0 22724 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_240
timestamp 1644511149
transform 1 0 23184 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_245
timestamp 1644511149
transform 1 0 23644 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_250
timestamp 1644511149
transform 1 0 24104 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_269
timestamp 1644511149
transform 1 0 25852 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_287
timestamp 1644511149
transform 1 0 27508 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1644511149
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1644511149
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_27
timestamp 1644511149
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_39
timestamp 1644511149
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1644511149
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1644511149
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_57
timestamp 1644511149
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_69
timestamp 1644511149
transform 1 0 7452 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_89
timestamp 1644511149
transform 1 0 9292 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_107
timestamp 1644511149
transform 1 0 10948 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1644511149
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_113
timestamp 1644511149
transform 1 0 11500 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_119
timestamp 1644511149
transform 1 0 12052 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_125
timestamp 1644511149
transform 1 0 12604 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_129
timestamp 1644511149
transform 1 0 12972 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_133
timestamp 1644511149
transform 1 0 13340 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_138
timestamp 1644511149
transform 1 0 13800 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_142
timestamp 1644511149
transform 1 0 14168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_145
timestamp 1644511149
transform 1 0 14444 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_149
timestamp 1644511149
transform 1 0 14812 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_159
timestamp 1644511149
transform 1 0 15732 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_166
timestamp 1644511149
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_179
timestamp 1644511149
transform 1 0 17572 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_187
timestamp 1644511149
transform 1 0 18308 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_191
timestamp 1644511149
transform 1 0 18676 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_202
timestamp 1644511149
transform 1 0 19688 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_209
timestamp 1644511149
transform 1 0 20332 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_216
timestamp 1644511149
transform 1 0 20976 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_222
timestamp 1644511149
transform 1 0 21528 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_228
timestamp 1644511149
transform 1 0 22080 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_240
timestamp 1644511149
transform 1 0 23184 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_247
timestamp 1644511149
transform 1 0 23828 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_251
timestamp 1644511149
transform 1 0 24196 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_255
timestamp 1644511149
transform 1 0 24564 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_259
timestamp 1644511149
transform 1 0 24932 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_263
timestamp 1644511149
transform 1 0 25300 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_275
timestamp 1644511149
transform 1 0 26404 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 1644511149
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_281
timestamp 1644511149
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_293
timestamp 1644511149
transform 1 0 28060 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1644511149
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1644511149
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1644511149
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_29
timestamp 1644511149
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_41
timestamp 1644511149
transform 1 0 4876 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_47
timestamp 1644511149
transform 1 0 5428 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_65
timestamp 1644511149
transform 1 0 7084 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_76
timestamp 1644511149
transform 1 0 8096 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_81
timestamp 1644511149
transform 1 0 8556 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_24_85
timestamp 1644511149
transform 1 0 8924 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_24_94
timestamp 1644511149
transform 1 0 9752 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_106
timestamp 1644511149
transform 1 0 10856 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_113
timestamp 1644511149
transform 1 0 11500 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_131
timestamp 1644511149
transform 1 0 13156 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_138
timestamp 1644511149
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_158
timestamp 1644511149
transform 1 0 15640 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_180
timestamp 1644511149
transform 1 0 17664 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_192
timestamp 1644511149
transform 1 0 18768 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_207
timestamp 1644511149
transform 1 0 20148 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_215
timestamp 1644511149
transform 1 0 20884 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_222
timestamp 1644511149
transform 1 0 21528 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_229
timestamp 1644511149
transform 1 0 22172 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_236
timestamp 1644511149
transform 1 0 22816 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_246
timestamp 1644511149
transform 1 0 23736 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_250
timestamp 1644511149
transform 1 0 24104 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_269
timestamp 1644511149
transform 1 0 25852 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_281
timestamp 1644511149
transform 1 0 26956 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_293
timestamp 1644511149
transform 1 0 28060 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_297
timestamp 1644511149
transform 1 0 28428 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1644511149
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_15
timestamp 1644511149
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_27
timestamp 1644511149
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_39
timestamp 1644511149
transform 1 0 4692 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_47
timestamp 1644511149
transform 1 0 5428 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_54
timestamp 1644511149
transform 1 0 6072 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_57
timestamp 1644511149
transform 1 0 6348 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_65
timestamp 1644511149
transform 1 0 7084 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_76
timestamp 1644511149
transform 1 0 8096 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_25_87
timestamp 1644511149
transform 1 0 9108 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_105
timestamp 1644511149
transform 1 0 10764 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_110
timestamp 1644511149
transform 1 0 11224 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_122
timestamp 1644511149
transform 1 0 12328 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_130
timestamp 1644511149
transform 1 0 13064 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_137
timestamp 1644511149
transform 1 0 13708 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_147
timestamp 1644511149
transform 1 0 14628 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_156
timestamp 1644511149
transform 1 0 15456 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_166
timestamp 1644511149
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_171
timestamp 1644511149
transform 1 0 16836 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_183
timestamp 1644511149
transform 1 0 17940 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_189
timestamp 1644511149
transform 1 0 18492 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_201
timestamp 1644511149
transform 1 0 19596 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_209
timestamp 1644511149
transform 1 0 20332 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_220
timestamp 1644511149
transform 1 0 21344 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_233
timestamp 1644511149
transform 1 0 22540 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_237
timestamp 1644511149
transform 1 0 22908 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_246
timestamp 1644511149
transform 1 0 23736 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_264
timestamp 1644511149
transform 1 0 25392 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_268
timestamp 1644511149
transform 1 0 25760 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_281
timestamp 1644511149
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_293
timestamp 1644511149
transform 1 0 28060 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_26_7
timestamp 1644511149
transform 1 0 1748 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_19
timestamp 1644511149
transform 1 0 2852 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1644511149
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_29
timestamp 1644511149
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_41
timestamp 1644511149
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_53
timestamp 1644511149
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_65
timestamp 1644511149
transform 1 0 7084 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_82
timestamp 1644511149
transform 1 0 8648 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_85
timestamp 1644511149
transform 1 0 8924 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_97
timestamp 1644511149
transform 1 0 10028 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_106
timestamp 1644511149
transform 1 0 10856 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_112
timestamp 1644511149
transform 1 0 11408 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_118
timestamp 1644511149
transform 1 0 11960 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_122
timestamp 1644511149
transform 1 0 12328 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_130
timestamp 1644511149
transform 1 0 13064 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_138
timestamp 1644511149
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_148
timestamp 1644511149
transform 1 0 14720 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_156
timestamp 1644511149
transform 1 0 15456 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_165
timestamp 1644511149
transform 1 0 16284 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_169
timestamp 1644511149
transform 1 0 16652 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_177
timestamp 1644511149
transform 1 0 17388 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_188
timestamp 1644511149
transform 1 0 18400 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_194
timestamp 1644511149
transform 1 0 18952 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_204
timestamp 1644511149
transform 1 0 19872 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_208
timestamp 1644511149
transform 1 0 20240 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_214
timestamp 1644511149
transform 1 0 20792 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_221
timestamp 1644511149
transform 1 0 21436 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_232
timestamp 1644511149
transform 1 0 22448 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_238
timestamp 1644511149
transform 1 0 23000 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_248
timestamp 1644511149
transform 1 0 23920 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_258
timestamp 1644511149
transform 1 0 24840 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_262
timestamp 1644511149
transform 1 0 25208 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_274
timestamp 1644511149
transform 1 0 26312 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_286
timestamp 1644511149
transform 1 0 27416 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_297
timestamp 1644511149
transform 1 0 28428 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_6
timestamp 1644511149
transform 1 0 1656 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_18
timestamp 1644511149
transform 1 0 2760 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_30
timestamp 1644511149
transform 1 0 3864 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_42
timestamp 1644511149
transform 1 0 4968 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_50
timestamp 1644511149
transform 1 0 5704 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_54
timestamp 1644511149
transform 1 0 6072 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_62
timestamp 1644511149
transform 1 0 6808 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_73
timestamp 1644511149
transform 1 0 7820 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_79
timestamp 1644511149
transform 1 0 8372 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_83
timestamp 1644511149
transform 1 0 8740 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_90
timestamp 1644511149
transform 1 0 9384 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_27_97
timestamp 1644511149
transform 1 0 10028 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_27_109
timestamp 1644511149
transform 1 0 11132 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_129
timestamp 1644511149
transform 1 0 12972 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_135
timestamp 1644511149
transform 1 0 13524 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_146
timestamp 1644511149
transform 1 0 14536 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_153
timestamp 1644511149
transform 1 0 15180 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_165
timestamp 1644511149
transform 1 0 16284 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_169
timestamp 1644511149
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_173
timestamp 1644511149
transform 1 0 17020 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_184
timestamp 1644511149
transform 1 0 18032 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_192
timestamp 1644511149
transform 1 0 18768 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_196
timestamp 1644511149
transform 1 0 19136 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_200
timestamp 1644511149
transform 1 0 19504 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_217
timestamp 1644511149
transform 1 0 21068 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_222
timestamp 1644511149
transform 1 0 21528 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_230
timestamp 1644511149
transform 1 0 22264 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_244
timestamp 1644511149
transform 1 0 23552 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_264
timestamp 1644511149
transform 1 0 25392 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_276
timestamp 1644511149
transform 1 0 26496 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_281
timestamp 1644511149
transform 1 0 26956 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_291
timestamp 1644511149
transform 1 0 27876 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_297
timestamp 1644511149
transform 1 0 28428 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_3
timestamp 1644511149
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_15
timestamp 1644511149
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1644511149
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_29
timestamp 1644511149
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_41
timestamp 1644511149
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_69
timestamp 1644511149
transform 1 0 7452 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_73
timestamp 1644511149
transform 1 0 7820 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_78
timestamp 1644511149
transform 1 0 8280 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_28_101
timestamp 1644511149
transform 1 0 10396 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_105
timestamp 1644511149
transform 1 0 10764 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_110
timestamp 1644511149
transform 1 0 11224 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_114
timestamp 1644511149
transform 1 0 11592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_118
timestamp 1644511149
transform 1 0 11960 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_123
timestamp 1644511149
transform 1 0 12420 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_130
timestamp 1644511149
transform 1 0 13064 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_137
timestamp 1644511149
transform 1 0 13708 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_149
timestamp 1644511149
transform 1 0 14812 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_153
timestamp 1644511149
transform 1 0 15180 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_162
timestamp 1644511149
transform 1 0 16008 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_166
timestamp 1644511149
transform 1 0 16376 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_184
timestamp 1644511149
transform 1 0 18032 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_28_193
timestamp 1644511149
transform 1 0 18860 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_206
timestamp 1644511149
transform 1 0 20056 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_216
timestamp 1644511149
transform 1 0 20976 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_220
timestamp 1644511149
transform 1 0 21344 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_228
timestamp 1644511149
transform 1 0 22080 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_234
timestamp 1644511149
transform 1 0 22632 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_242
timestamp 1644511149
transform 1 0 23368 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_249
timestamp 1644511149
transform 1 0 24012 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_255
timestamp 1644511149
transform 1 0 24564 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_267
timestamp 1644511149
transform 1 0 25668 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_279
timestamp 1644511149
transform 1 0 26772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_291
timestamp 1644511149
transform 1 0 27876 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1644511149
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_15
timestamp 1644511149
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_27
timestamp 1644511149
transform 1 0 3588 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_35
timestamp 1644511149
transform 1 0 4324 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_54
timestamp 1644511149
transform 1 0 6072 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_57
timestamp 1644511149
transform 1 0 6348 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_29_66
timestamp 1644511149
transform 1 0 7176 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_78
timestamp 1644511149
transform 1 0 8280 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_84
timestamp 1644511149
transform 1 0 8832 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_96
timestamp 1644511149
transform 1 0 9936 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_100
timestamp 1644511149
transform 1 0 10304 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_106
timestamp 1644511149
transform 1 0 10856 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_29_129
timestamp 1644511149
transform 1 0 12972 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_136
timestamp 1644511149
transform 1 0 13616 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_145
timestamp 1644511149
transform 1 0 14444 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_154
timestamp 1644511149
transform 1 0 15272 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_166
timestamp 1644511149
transform 1 0 16376 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_179
timestamp 1644511149
transform 1 0 17572 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_183
timestamp 1644511149
transform 1 0 17940 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_202
timestamp 1644511149
transform 1 0 19688 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_206
timestamp 1644511149
transform 1 0 20056 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_213
timestamp 1644511149
transform 1 0 20700 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_220
timestamp 1644511149
transform 1 0 21344 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_29_233
timestamp 1644511149
transform 1 0 22540 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_244
timestamp 1644511149
transform 1 0 23552 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_262
timestamp 1644511149
transform 1 0 25208 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_274
timestamp 1644511149
transform 1 0 26312 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_29_281
timestamp 1644511149
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_293
timestamp 1644511149
transform 1 0 28060 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_30_6
timestamp 1644511149
transform 1 0 1656 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_18
timestamp 1644511149
transform 1 0 2760 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_26
timestamp 1644511149
transform 1 0 3496 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_29
timestamp 1644511149
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_41
timestamp 1644511149
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_53
timestamp 1644511149
transform 1 0 5980 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_59
timestamp 1644511149
transform 1 0 6532 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_76
timestamp 1644511149
transform 1 0 8096 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_30_94
timestamp 1644511149
transform 1 0 9752 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_100
timestamp 1644511149
transform 1 0 10304 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_110
timestamp 1644511149
transform 1 0 11224 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_115
timestamp 1644511149
transform 1 0 11684 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_30_126
timestamp 1644511149
transform 1 0 12696 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1644511149
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1644511149
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_149
timestamp 1644511149
transform 1 0 14812 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_158
timestamp 1644511149
transform 1 0 15640 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_167
timestamp 1644511149
transform 1 0 16468 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_173
timestamp 1644511149
transform 1 0 17020 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_183
timestamp 1644511149
transform 1 0 17940 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_188
timestamp 1644511149
transform 1 0 18400 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_194
timestamp 1644511149
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_197
timestamp 1644511149
transform 1 0 19228 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_204
timestamp 1644511149
transform 1 0 19872 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_214
timestamp 1644511149
transform 1 0 20792 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_218
timestamp 1644511149
transform 1 0 21160 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_227
timestamp 1644511149
transform 1 0 21988 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_234
timestamp 1644511149
transform 1 0 22632 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_238
timestamp 1644511149
transform 1 0 23000 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_248
timestamp 1644511149
transform 1 0 23920 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_269
timestamp 1644511149
transform 1 0 25852 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_281
timestamp 1644511149
transform 1 0 26956 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_293
timestamp 1644511149
transform 1 0 28060 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_31_5
timestamp 1644511149
transform 1 0 1564 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_17
timestamp 1644511149
transform 1 0 2668 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_29
timestamp 1644511149
transform 1 0 3772 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_41
timestamp 1644511149
transform 1 0 4876 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_53
timestamp 1644511149
transform 1 0 5980 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_57
timestamp 1644511149
transform 1 0 6348 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_61
timestamp 1644511149
transform 1 0 6716 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_65
timestamp 1644511149
transform 1 0 7084 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_31_73
timestamp 1644511149
transform 1 0 7820 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_81
timestamp 1644511149
transform 1 0 8556 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_87
timestamp 1644511149
transform 1 0 9108 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_92
timestamp 1644511149
transform 1 0 9568 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_96
timestamp 1644511149
transform 1 0 9936 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_100
timestamp 1644511149
transform 1 0 10304 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_110
timestamp 1644511149
transform 1 0 11224 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_116
timestamp 1644511149
transform 1 0 11776 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_130
timestamp 1644511149
transform 1 0 13064 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_137
timestamp 1644511149
transform 1 0 13708 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_145
timestamp 1644511149
transform 1 0 14444 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_150
timestamp 1644511149
transform 1 0 14904 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_158
timestamp 1644511149
transform 1 0 15640 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_166
timestamp 1644511149
transform 1 0 16376 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_175
timestamp 1644511149
transform 1 0 17204 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_31_194
timestamp 1644511149
transform 1 0 18952 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_213
timestamp 1644511149
transform 1 0 20700 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_222
timestamp 1644511149
transform 1 0 21528 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_225
timestamp 1644511149
transform 1 0 21804 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_234
timestamp 1644511149
transform 1 0 22632 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_241
timestamp 1644511149
transform 1 0 23276 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_248
timestamp 1644511149
transform 1 0 23920 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_254
timestamp 1644511149
transform 1 0 24472 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_258
timestamp 1644511149
transform 1 0 24840 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_270
timestamp 1644511149
transform 1 0 25944 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_278
timestamp 1644511149
transform 1 0 26680 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_281
timestamp 1644511149
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_293
timestamp 1644511149
transform 1 0 28060 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_13
timestamp 1644511149
transform 1 0 2300 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_25
timestamp 1644511149
transform 1 0 3404 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_29
timestamp 1644511149
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_41
timestamp 1644511149
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_53
timestamp 1644511149
transform 1 0 5980 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_64
timestamp 1644511149
transform 1 0 6992 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_71
timestamp 1644511149
transform 1 0 7636 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_82
timestamp 1644511149
transform 1 0 8648 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_85
timestamp 1644511149
transform 1 0 8924 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_102
timestamp 1644511149
transform 1 0 10488 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_106
timestamp 1644511149
transform 1 0 10856 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_123
timestamp 1644511149
transform 1 0 12420 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_127
timestamp 1644511149
transform 1 0 12788 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_138
timestamp 1644511149
transform 1 0 13800 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_157
timestamp 1644511149
transform 1 0 15548 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_165
timestamp 1644511149
transform 1 0 16284 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_179
timestamp 1644511149
transform 1 0 17572 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_191
timestamp 1644511149
transform 1 0 18676 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1644511149
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_199
timestamp 1644511149
transform 1 0 19412 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_204
timestamp 1644511149
transform 1 0 19872 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_208
timestamp 1644511149
transform 1 0 20240 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_212
timestamp 1644511149
transform 1 0 20608 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_216
timestamp 1644511149
transform 1 0 20976 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_219
timestamp 1644511149
transform 1 0 21252 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_225
timestamp 1644511149
transform 1 0 21804 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_229
timestamp 1644511149
transform 1 0 22172 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_247
timestamp 1644511149
transform 1 0 23828 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1644511149
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_253
timestamp 1644511149
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_265
timestamp 1644511149
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_277
timestamp 1644511149
transform 1 0 26588 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_289
timestamp 1644511149
transform 1 0 27692 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_297
timestamp 1644511149
transform 1 0 28428 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1644511149
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_15
timestamp 1644511149
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_27
timestamp 1644511149
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_39
timestamp 1644511149
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1644511149
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1644511149
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_57
timestamp 1644511149
transform 1 0 6348 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_61
timestamp 1644511149
transform 1 0 6716 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_78
timestamp 1644511149
transform 1 0 8280 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_82
timestamp 1644511149
transform 1 0 8648 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_87
timestamp 1644511149
transform 1 0 9108 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_94
timestamp 1644511149
transform 1 0 9752 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_103
timestamp 1644511149
transform 1 0 10580 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_110
timestamp 1644511149
transform 1 0 11224 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_113
timestamp 1644511149
transform 1 0 11500 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_33_125
timestamp 1644511149
transform 1 0 12604 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_33_135
timestamp 1644511149
transform 1 0 13524 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_140
timestamp 1644511149
transform 1 0 13984 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_144
timestamp 1644511149
transform 1 0 14352 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_155
timestamp 1644511149
transform 1 0 15364 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_161
timestamp 1644511149
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1644511149
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_185
timestamp 1644511149
transform 1 0 18124 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_197
timestamp 1644511149
transform 1 0 19228 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_202
timestamp 1644511149
transform 1 0 19688 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_213
timestamp 1644511149
transform 1 0 20700 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_218
timestamp 1644511149
transform 1 0 21160 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_33_241
timestamp 1644511149
transform 1 0 23276 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_253
timestamp 1644511149
transform 1 0 24380 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_265
timestamp 1644511149
transform 1 0 25484 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_277
timestamp 1644511149
transform 1 0 26588 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_281
timestamp 1644511149
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_293
timestamp 1644511149
transform 1 0 28060 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1644511149
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1644511149
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1644511149
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_29
timestamp 1644511149
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_41
timestamp 1644511149
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_53
timestamp 1644511149
transform 1 0 5980 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_61
timestamp 1644511149
transform 1 0 6716 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_64
timestamp 1644511149
transform 1 0 6992 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_71
timestamp 1644511149
transform 1 0 7636 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_82
timestamp 1644511149
transform 1 0 8648 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_85
timestamp 1644511149
transform 1 0 8924 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_89
timestamp 1644511149
transform 1 0 9292 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_99
timestamp 1644511149
transform 1 0 10212 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_103
timestamp 1644511149
transform 1 0 10580 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_110
timestamp 1644511149
transform 1 0 11224 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_115
timestamp 1644511149
transform 1 0 11684 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 1644511149
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1644511149
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_143
timestamp 1644511149
transform 1 0 14260 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_155
timestamp 1644511149
transform 1 0 15364 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_161
timestamp 1644511149
transform 1 0 15916 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_172
timestamp 1644511149
transform 1 0 16928 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_179
timestamp 1644511149
transform 1 0 17572 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_183
timestamp 1644511149
transform 1 0 17940 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_194
timestamp 1644511149
transform 1 0 18952 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_197
timestamp 1644511149
transform 1 0 19228 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_203
timestamp 1644511149
transform 1 0 19780 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_214
timestamp 1644511149
transform 1 0 20792 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_232
timestamp 1644511149
transform 1 0 22448 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_250
timestamp 1644511149
transform 1 0 24104 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_253
timestamp 1644511149
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_265
timestamp 1644511149
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_277
timestamp 1644511149
transform 1 0 26588 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_289
timestamp 1644511149
transform 1 0 27692 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_297
timestamp 1644511149
transform 1 0 28428 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_6
timestamp 1644511149
transform 1 0 1656 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_18
timestamp 1644511149
transform 1 0 2760 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_30
timestamp 1644511149
transform 1 0 3864 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_42
timestamp 1644511149
transform 1 0 4968 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_54
timestamp 1644511149
transform 1 0 6072 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_57
timestamp 1644511149
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_69
timestamp 1644511149
transform 1 0 7452 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_87
timestamp 1644511149
transform 1 0 9108 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_105
timestamp 1644511149
transform 1 0 10764 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_110
timestamp 1644511149
transform 1 0 11224 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_122
timestamp 1644511149
transform 1 0 12328 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_129
timestamp 1644511149
transform 1 0 12972 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_133
timestamp 1644511149
transform 1 0 13340 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_144
timestamp 1644511149
transform 1 0 14352 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_157
timestamp 1644511149
transform 1 0 15548 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_164
timestamp 1644511149
transform 1 0 16192 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_172
timestamp 1644511149
transform 1 0 16928 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_176
timestamp 1644511149
transform 1 0 17296 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_194
timestamp 1644511149
transform 1 0 18952 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_201
timestamp 1644511149
transform 1 0 19596 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_210
timestamp 1644511149
transform 1 0 20424 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_214
timestamp 1644511149
transform 1 0 20792 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_218
timestamp 1644511149
transform 1 0 21160 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_222
timestamp 1644511149
transform 1 0 21528 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_225
timestamp 1644511149
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_237
timestamp 1644511149
transform 1 0 22908 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_249
timestamp 1644511149
transform 1 0 24012 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_261
timestamp 1644511149
transform 1 0 25116 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_273
timestamp 1644511149
transform 1 0 26220 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1644511149
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_281
timestamp 1644511149
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_293
timestamp 1644511149
transform 1 0 28060 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_36_3
timestamp 1644511149
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_15
timestamp 1644511149
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1644511149
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_29
timestamp 1644511149
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_41
timestamp 1644511149
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_53
timestamp 1644511149
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_65
timestamp 1644511149
transform 1 0 7084 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_36_76
timestamp 1644511149
transform 1 0 8096 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_85
timestamp 1644511149
transform 1 0 8924 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_89
timestamp 1644511149
transform 1 0 9292 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_93
timestamp 1644511149
transform 1 0 9660 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_97
timestamp 1644511149
transform 1 0 10028 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_102
timestamp 1644511149
transform 1 0 10488 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_120
timestamp 1644511149
transform 1 0 12144 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_138
timestamp 1644511149
transform 1 0 13800 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_141
timestamp 1644511149
transform 1 0 14076 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_159
timestamp 1644511149
transform 1 0 15732 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_163
timestamp 1644511149
transform 1 0 16100 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_36_173
timestamp 1644511149
transform 1 0 17020 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_184
timestamp 1644511149
transform 1 0 18032 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_188
timestamp 1644511149
transform 1 0 18400 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_194
timestamp 1644511149
transform 1 0 18952 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_206
timestamp 1644511149
transform 1 0 20056 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_217
timestamp 1644511149
transform 1 0 21068 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_222
timestamp 1644511149
transform 1 0 21528 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_226
timestamp 1644511149
transform 1 0 21896 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_238
timestamp 1644511149
transform 1 0 23000 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_250
timestamp 1644511149
transform 1 0 24104 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_253
timestamp 1644511149
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_265
timestamp 1644511149
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_277
timestamp 1644511149
transform 1 0 26588 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_289
timestamp 1644511149
transform 1 0 27692 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_297
timestamp 1644511149
transform 1 0 28428 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_3
timestamp 1644511149
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_15
timestamp 1644511149
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_27
timestamp 1644511149
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_39
timestamp 1644511149
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1644511149
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1644511149
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_57
timestamp 1644511149
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_69
timestamp 1644511149
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_81
timestamp 1644511149
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_93
timestamp 1644511149
transform 1 0 9660 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_101
timestamp 1644511149
transform 1 0 10396 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_104
timestamp 1644511149
transform 1 0 10672 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_37_113
timestamp 1644511149
transform 1 0 11500 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_126
timestamp 1644511149
transform 1 0 12696 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_144
timestamp 1644511149
transform 1 0 14352 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_155
timestamp 1644511149
transform 1 0 15364 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_164
timestamp 1644511149
transform 1 0 16192 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_185
timestamp 1644511149
transform 1 0 18124 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_203
timestamp 1644511149
transform 1 0 19780 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_222
timestamp 1644511149
transform 1 0 21528 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_225
timestamp 1644511149
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_237
timestamp 1644511149
transform 1 0 22908 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_249
timestamp 1644511149
transform 1 0 24012 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_261
timestamp 1644511149
transform 1 0 25116 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_273
timestamp 1644511149
transform 1 0 26220 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1644511149
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_281
timestamp 1644511149
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_293
timestamp 1644511149
transform 1 0 28060 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_38_3
timestamp 1644511149
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_15
timestamp 1644511149
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1644511149
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_29
timestamp 1644511149
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_41
timestamp 1644511149
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_53
timestamp 1644511149
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_65
timestamp 1644511149
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1644511149
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1644511149
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_85
timestamp 1644511149
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_97
timestamp 1644511149
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_109
timestamp 1644511149
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_121
timestamp 1644511149
transform 1 0 12236 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_38_130
timestamp 1644511149
transform 1 0 13064 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_135
timestamp 1644511149
transform 1 0 13524 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1644511149
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_141
timestamp 1644511149
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_155
timestamp 1644511149
transform 1 0 15364 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_162
timestamp 1644511149
transform 1 0 16008 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_173
timestamp 1644511149
transform 1 0 17020 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_179
timestamp 1644511149
transform 1 0 17572 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_184
timestamp 1644511149
transform 1 0 18032 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_189
timestamp 1644511149
transform 1 0 18492 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_194
timestamp 1644511149
transform 1 0 18952 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_197
timestamp 1644511149
transform 1 0 19228 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_203
timestamp 1644511149
transform 1 0 19780 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_211
timestamp 1644511149
transform 1 0 20516 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_223
timestamp 1644511149
transform 1 0 21620 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_235
timestamp 1644511149
transform 1 0 22724 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_247
timestamp 1644511149
transform 1 0 23828 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp 1644511149
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_253
timestamp 1644511149
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_265
timestamp 1644511149
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_277
timestamp 1644511149
transform 1 0 26588 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_289
timestamp 1644511149
transform 1 0 27692 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_297
timestamp 1644511149
transform 1 0 28428 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_6
timestamp 1644511149
transform 1 0 1656 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_18
timestamp 1644511149
transform 1 0 2760 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_30
timestamp 1644511149
transform 1 0 3864 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_42
timestamp 1644511149
transform 1 0 4968 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_54
timestamp 1644511149
transform 1 0 6072 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_57
timestamp 1644511149
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_69
timestamp 1644511149
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_81
timestamp 1644511149
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_93
timestamp 1644511149
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1644511149
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1644511149
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_113
timestamp 1644511149
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_125
timestamp 1644511149
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_137
timestamp 1644511149
transform 1 0 13708 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_39_148
timestamp 1644511149
transform 1 0 14720 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_159
timestamp 1644511149
transform 1 0 15732 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_166
timestamp 1644511149
transform 1 0 16376 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_185
timestamp 1644511149
transform 1 0 18124 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_197
timestamp 1644511149
transform 1 0 19228 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_202
timestamp 1644511149
transform 1 0 19688 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_39_206
timestamp 1644511149
transform 1 0 20056 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_39_216
timestamp 1644511149
transform 1 0 20976 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_39_225
timestamp 1644511149
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_237
timestamp 1644511149
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_249
timestamp 1644511149
transform 1 0 24012 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_261
timestamp 1644511149
transform 1 0 25116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_273
timestamp 1644511149
transform 1 0 26220 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1644511149
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_281
timestamp 1644511149
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_293
timestamp 1644511149
transform 1 0 28060 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_297
timestamp 1644511149
transform 1 0 28428 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_40_3
timestamp 1644511149
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_15
timestamp 1644511149
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1644511149
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_29
timestamp 1644511149
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_41
timestamp 1644511149
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_53
timestamp 1644511149
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_65
timestamp 1644511149
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1644511149
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1644511149
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_85
timestamp 1644511149
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_97
timestamp 1644511149
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_109
timestamp 1644511149
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_121
timestamp 1644511149
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 1644511149
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1644511149
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_40_141
timestamp 1644511149
transform 1 0 14076 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_160
timestamp 1644511149
transform 1 0 15824 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_164
timestamp 1644511149
transform 1 0 16192 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_168
timestamp 1644511149
transform 1 0 16560 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_172
timestamp 1644511149
transform 1 0 16928 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_40_176
timestamp 1644511149
transform 1 0 17296 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_188
timestamp 1644511149
transform 1 0 18400 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_197
timestamp 1644511149
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_209
timestamp 1644511149
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_221
timestamp 1644511149
transform 1 0 21436 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_233
timestamp 1644511149
transform 1 0 22540 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_245
timestamp 1644511149
transform 1 0 23644 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1644511149
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_253
timestamp 1644511149
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_265
timestamp 1644511149
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_277
timestamp 1644511149
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_289
timestamp 1644511149
transform 1 0 27692 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_297
timestamp 1644511149
transform 1 0 28428 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_7
timestamp 1644511149
transform 1 0 1748 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_11
timestamp 1644511149
transform 1 0 2116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_23
timestamp 1644511149
transform 1 0 3220 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_35
timestamp 1644511149
transform 1 0 4324 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_47
timestamp 1644511149
transform 1 0 5428 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1644511149
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_57
timestamp 1644511149
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_69
timestamp 1644511149
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_81
timestamp 1644511149
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_93
timestamp 1644511149
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1644511149
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1644511149
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_113
timestamp 1644511149
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_125
timestamp 1644511149
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_137
timestamp 1644511149
transform 1 0 13708 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_145
timestamp 1644511149
transform 1 0 14444 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_151
timestamp 1644511149
transform 1 0 14996 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_163
timestamp 1644511149
transform 1 0 16100 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1644511149
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_169
timestamp 1644511149
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_181
timestamp 1644511149
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_193
timestamp 1644511149
transform 1 0 18860 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_205
timestamp 1644511149
transform 1 0 19964 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_217
timestamp 1644511149
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 1644511149
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_225
timestamp 1644511149
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_237
timestamp 1644511149
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_249
timestamp 1644511149
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_261
timestamp 1644511149
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_273
timestamp 1644511149
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1644511149
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_281
timestamp 1644511149
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_293
timestamp 1644511149
transform 1 0 28060 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_3
timestamp 1644511149
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_15
timestamp 1644511149
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1644511149
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_29
timestamp 1644511149
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_41
timestamp 1644511149
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_53
timestamp 1644511149
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_65
timestamp 1644511149
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1644511149
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1644511149
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_85
timestamp 1644511149
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_97
timestamp 1644511149
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_109
timestamp 1644511149
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_121
timestamp 1644511149
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_133
timestamp 1644511149
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1644511149
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_141
timestamp 1644511149
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_153
timestamp 1644511149
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_165
timestamp 1644511149
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_177
timestamp 1644511149
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_189
timestamp 1644511149
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1644511149
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_197
timestamp 1644511149
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_209
timestamp 1644511149
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_221
timestamp 1644511149
transform 1 0 21436 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_233
timestamp 1644511149
transform 1 0 22540 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_245
timestamp 1644511149
transform 1 0 23644 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1644511149
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_253
timestamp 1644511149
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_265
timestamp 1644511149
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_277
timestamp 1644511149
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_291
timestamp 1644511149
transform 1 0 27876 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_297
timestamp 1644511149
transform 1 0 28428 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_43_3
timestamp 1644511149
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_15
timestamp 1644511149
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_27
timestamp 1644511149
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_39
timestamp 1644511149
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1644511149
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1644511149
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_57
timestamp 1644511149
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_69
timestamp 1644511149
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_81
timestamp 1644511149
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_93
timestamp 1644511149
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1644511149
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1644511149
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_113
timestamp 1644511149
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_125
timestamp 1644511149
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_137
timestamp 1644511149
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_149
timestamp 1644511149
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_161
timestamp 1644511149
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1644511149
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_169
timestamp 1644511149
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_181
timestamp 1644511149
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_193
timestamp 1644511149
transform 1 0 18860 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_205
timestamp 1644511149
transform 1 0 19964 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_217
timestamp 1644511149
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1644511149
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_225
timestamp 1644511149
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_237
timestamp 1644511149
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_249
timestamp 1644511149
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_261
timestamp 1644511149
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_273
timestamp 1644511149
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1644511149
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_281
timestamp 1644511149
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_293
timestamp 1644511149
transform 1 0 28060 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_44_6
timestamp 1644511149
transform 1 0 1656 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_18
timestamp 1644511149
transform 1 0 2760 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_26
timestamp 1644511149
transform 1 0 3496 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_44_29
timestamp 1644511149
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_41
timestamp 1644511149
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_53
timestamp 1644511149
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_65
timestamp 1644511149
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1644511149
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1644511149
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_85
timestamp 1644511149
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_97
timestamp 1644511149
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_109
timestamp 1644511149
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_121
timestamp 1644511149
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 1644511149
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1644511149
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_141
timestamp 1644511149
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_153
timestamp 1644511149
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_165
timestamp 1644511149
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_177
timestamp 1644511149
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_189
timestamp 1644511149
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1644511149
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_197
timestamp 1644511149
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_209
timestamp 1644511149
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_221
timestamp 1644511149
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_233
timestamp 1644511149
transform 1 0 22540 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_245
timestamp 1644511149
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1644511149
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_253
timestamp 1644511149
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_265
timestamp 1644511149
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_277
timestamp 1644511149
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_289
timestamp 1644511149
transform 1 0 27692 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_293
timestamp 1644511149
transform 1 0 28060 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_297
timestamp 1644511149
transform 1 0 28428 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_7
timestamp 1644511149
transform 1 0 1748 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_11
timestamp 1644511149
transform 1 0 2116 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_45_15
timestamp 1644511149
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_27
timestamp 1644511149
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_39
timestamp 1644511149
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1644511149
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1644511149
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_57
timestamp 1644511149
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_69
timestamp 1644511149
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_81
timestamp 1644511149
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_93
timestamp 1644511149
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 1644511149
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1644511149
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_113
timestamp 1644511149
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_125
timestamp 1644511149
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_137
timestamp 1644511149
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_149
timestamp 1644511149
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_161
timestamp 1644511149
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1644511149
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_169
timestamp 1644511149
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_181
timestamp 1644511149
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_193
timestamp 1644511149
transform 1 0 18860 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_205
timestamp 1644511149
transform 1 0 19964 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_217
timestamp 1644511149
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1644511149
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_45_225
timestamp 1644511149
transform 1 0 21804 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_45_244
timestamp 1644511149
transform 1 0 23552 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_45_262
timestamp 1644511149
transform 1 0 25208 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_274
timestamp 1644511149
transform 1 0 26312 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_45_281
timestamp 1644511149
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_297
timestamp 1644511149
transform 1 0 28428 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_3
timestamp 1644511149
transform 1 0 1380 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_11
timestamp 1644511149
transform 1 0 2116 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_15
timestamp 1644511149
transform 1 0 2484 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_23
timestamp 1644511149
transform 1 0 3220 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1644511149
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_29
timestamp 1644511149
transform 1 0 3772 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_46_34
timestamp 1644511149
transform 1 0 4232 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_46
timestamp 1644511149
transform 1 0 5336 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_54
timestamp 1644511149
transform 1 0 6072 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_46_57
timestamp 1644511149
transform 1 0 6348 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_69
timestamp 1644511149
transform 1 0 7452 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_81
timestamp 1644511149
transform 1 0 8556 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_85
timestamp 1644511149
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_97
timestamp 1644511149
transform 1 0 10028 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_105
timestamp 1644511149
transform 1 0 10764 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_46_109
timestamp 1644511149
transform 1 0 11132 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_113
timestamp 1644511149
transform 1 0 11500 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_125
timestamp 1644511149
transform 1 0 12604 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_137
timestamp 1644511149
transform 1 0 13708 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_141
timestamp 1644511149
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_153
timestamp 1644511149
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_165
timestamp 1644511149
transform 1 0 16284 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_173
timestamp 1644511149
transform 1 0 17020 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_185
timestamp 1644511149
transform 1 0 18124 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_193
timestamp 1644511149
transform 1 0 18860 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_46_197
timestamp 1644511149
transform 1 0 19228 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_46_202
timestamp 1644511149
transform 1 0 19688 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_214
timestamp 1644511149
transform 1 0 20792 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_222
timestamp 1644511149
transform 1 0 21528 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_228
timestamp 1644511149
transform 1 0 22080 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_232
timestamp 1644511149
transform 1 0 22448 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_240
timestamp 1644511149
transform 1 0 23184 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_250
timestamp 1644511149
transform 1 0 24104 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_253
timestamp 1644511149
transform 1 0 24380 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_261
timestamp 1644511149
transform 1 0 25116 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_267
timestamp 1644511149
transform 1 0 25668 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_272
timestamp 1644511149
transform 1 0 26128 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_46_281
timestamp 1644511149
transform 1 0 26956 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_287
timestamp 1644511149
transform 1 0 27508 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_291
timestamp 1644511149
transform 1 0 27876 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_297
timestamp 1644511149
transform 1 0 28428 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1644511149
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1644511149
transform -1 0 28888 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1644511149
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1644511149
transform -1 0 28888 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1644511149
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1644511149
transform -1 0 28888 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1644511149
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1644511149
transform -1 0 28888 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1644511149
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1644511149
transform -1 0 28888 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1644511149
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1644511149
transform -1 0 28888 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1644511149
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1644511149
transform -1 0 28888 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1644511149
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1644511149
transform -1 0 28888 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1644511149
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1644511149
transform -1 0 28888 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1644511149
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1644511149
transform -1 0 28888 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1644511149
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1644511149
transform -1 0 28888 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1644511149
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1644511149
transform -1 0 28888 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1644511149
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1644511149
transform -1 0 28888 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1644511149
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1644511149
transform -1 0 28888 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1644511149
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1644511149
transform -1 0 28888 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1644511149
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1644511149
transform -1 0 28888 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1644511149
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1644511149
transform -1 0 28888 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1644511149
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1644511149
transform -1 0 28888 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1644511149
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1644511149
transform -1 0 28888 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1644511149
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1644511149
transform -1 0 28888 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1644511149
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1644511149
transform -1 0 28888 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1644511149
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1644511149
transform -1 0 28888 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1644511149
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1644511149
transform -1 0 28888 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1644511149
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1644511149
transform -1 0 28888 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1644511149
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1644511149
transform -1 0 28888 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1644511149
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1644511149
transform -1 0 28888 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1644511149
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1644511149
transform -1 0 28888 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1644511149
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1644511149
transform -1 0 28888 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1644511149
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1644511149
transform -1 0 28888 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1644511149
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1644511149
transform -1 0 28888 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1644511149
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1644511149
transform -1 0 28888 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1644511149
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1644511149
transform -1 0 28888 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1644511149
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1644511149
transform -1 0 28888 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1644511149
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1644511149
transform -1 0 28888 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1644511149
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1644511149
transform -1 0 28888 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1644511149
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1644511149
transform -1 0 28888 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1644511149
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1644511149
transform -1 0 28888 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1644511149
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1644511149
transform -1 0 28888 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1644511149
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1644511149
transform -1 0 28888 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1644511149
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1644511149
transform -1 0 28888 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1644511149
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1644511149
transform -1 0 28888 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1644511149
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1644511149
transform -1 0 28888 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1644511149
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1644511149
transform -1 0 28888 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1644511149
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1644511149
transform -1 0 28888 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1644511149
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1644511149
transform -1 0 28888 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1644511149
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1644511149
transform -1 0 28888 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1644511149
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1644511149
transform -1 0 28888 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1644511149
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1644511149
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1644511149
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1644511149
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1644511149
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1644511149
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1644511149
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1644511149
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1644511149
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1644511149
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1644511149
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1644511149
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1644511149
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1644511149
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1644511149
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1644511149
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1644511149
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1644511149
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1644511149
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1644511149
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1644511149
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1644511149
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1644511149
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1644511149
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1644511149
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1644511149
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1644511149
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1644511149
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1644511149
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1644511149
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1644511149
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1644511149
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1644511149
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1644511149
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1644511149
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1644511149
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1644511149
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1644511149
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1644511149
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1644511149
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1644511149
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1644511149
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1644511149
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1644511149
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1644511149
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1644511149
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1644511149
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1644511149
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1644511149
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1644511149
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1644511149
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1644511149
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1644511149
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1644511149
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1644511149
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1644511149
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1644511149
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1644511149
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1644511149
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1644511149
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1644511149
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1644511149
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1644511149
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1644511149
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1644511149
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1644511149
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1644511149
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1644511149
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1644511149
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1644511149
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1644511149
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1644511149
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1644511149
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1644511149
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1644511149
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1644511149
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1644511149
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1644511149
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1644511149
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1644511149
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1644511149
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1644511149
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1644511149
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1644511149
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1644511149
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1644511149
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1644511149
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1644511149
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1644511149
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1644511149
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1644511149
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1644511149
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1644511149
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1644511149
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1644511149
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1644511149
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1644511149
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1644511149
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1644511149
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1644511149
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1644511149
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1644511149
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1644511149
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1644511149
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1644511149
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1644511149
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1644511149
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1644511149
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1644511149
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1644511149
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1644511149
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1644511149
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1644511149
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1644511149
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1644511149
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1644511149
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1644511149
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1644511149
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1644511149
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1644511149
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1644511149
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1644511149
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1644511149
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1644511149
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1644511149
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1644511149
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1644511149
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1644511149
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1644511149
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1644511149
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1644511149
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1644511149
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1644511149
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1644511149
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1644511149
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1644511149
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1644511149
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1644511149
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1644511149
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1644511149
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1644511149
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1644511149
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1644511149
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1644511149
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1644511149
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1644511149
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1644511149
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1644511149
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1644511149
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1644511149
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1644511149
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1644511149
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1644511149
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1644511149
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1644511149
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1644511149
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1644511149
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1644511149
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1644511149
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1644511149
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1644511149
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1644511149
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1644511149
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1644511149
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1644511149
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1644511149
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1644511149
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1644511149
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1644511149
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1644511149
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1644511149
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1644511149
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1644511149
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1644511149
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1644511149
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1644511149
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1644511149
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1644511149
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1644511149
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1644511149
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1644511149
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1644511149
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1644511149
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1644511149
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1644511149
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1644511149
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1644511149
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1644511149
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1644511149
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1644511149
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1644511149
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1644511149
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1644511149
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1644511149
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1644511149
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1644511149
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1644511149
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1644511149
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1644511149
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1644511149
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1644511149
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1644511149
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1644511149
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1644511149
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1644511149
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1644511149
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1644511149
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1644511149
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1644511149
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1644511149
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1644511149
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1644511149
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1644511149
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1644511149
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1644511149
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1644511149
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1644511149
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1644511149
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1644511149
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1644511149
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1644511149
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1644511149
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1644511149
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1644511149
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1644511149
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1644511149
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1644511149
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1644511149
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1644511149
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1644511149
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1644511149
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1644511149
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1644511149
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1644511149
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1644511149
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1644511149
transform 1 0 6256 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1644511149
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1644511149
transform 1 0 11408 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1644511149
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1644511149
transform 1 0 16560 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1644511149
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1644511149
transform 1 0 21712 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1644511149
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1644511149
transform 1 0 26864 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_1  _0524_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 15548 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0525_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17296 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0526_
timestamp 1644511149
transform 1 0 17940 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0527_
timestamp 1644511149
transform -1 0 19228 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__nor4_1  _0528_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20884 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0529_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19688 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0530_
timestamp 1644511149
transform 1 0 19044 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0531_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21896 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0532_
timestamp 1644511149
transform 1 0 22540 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__or4_2  _0533_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16836 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0534_
timestamp 1644511149
transform 1 0 17756 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _0535_
timestamp 1644511149
transform 1 0 18032 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0536_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 19504 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0537_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19688 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0538_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 20608 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0539_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22356 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__or3_1  _0540_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22448 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0541_
timestamp 1644511149
transform 1 0 24564 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0542_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 25576 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0543_
timestamp 1644511149
transform 1 0 25116 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0544_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25300 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0545_
timestamp 1644511149
transform -1 0 25668 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0546_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25852 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0547_
timestamp 1644511149
transform 1 0 24104 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0548_
timestamp 1644511149
transform 1 0 23644 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0549_
timestamp 1644511149
transform -1 0 23828 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0550_
timestamp 1644511149
transform 1 0 21160 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0551_
timestamp 1644511149
transform -1 0 25208 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0552_
timestamp 1644511149
transform 1 0 24656 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0553_
timestamp 1644511149
transform 1 0 23000 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0554_
timestamp 1644511149
transform -1 0 26220 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _0555_
timestamp 1644511149
transform 1 0 24656 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0556_
timestamp 1644511149
transform -1 0 26496 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0557_
timestamp 1644511149
transform 1 0 27232 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0558_
timestamp 1644511149
transform 1 0 25576 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0559_
timestamp 1644511149
transform -1 0 25576 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0560_
timestamp 1644511149
transform 1 0 26404 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0561_
timestamp 1644511149
transform 1 0 24104 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0562_
timestamp 1644511149
transform -1 0 23920 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0563_
timestamp 1644511149
transform 1 0 23828 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0564_
timestamp 1644511149
transform 1 0 21988 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0565_
timestamp 1644511149
transform -1 0 22448 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0566_
timestamp 1644511149
transform 1 0 22540 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0567_
timestamp 1644511149
transform 1 0 18308 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _0568_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17848 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__or3_2  _0569_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19228 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _0570_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 18400 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0571_
timestamp 1644511149
transform 1 0 19688 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0572_
timestamp 1644511149
transform -1 0 22908 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _0573_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 22172 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0574_
timestamp 1644511149
transform 1 0 7544 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__or4_2  _0575_
timestamp 1644511149
transform 1 0 10396 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or4_2  _0576_
timestamp 1644511149
transform -1 0 13708 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nor4_4  _0577_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 10120 0 1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__or3_1  _0578_
timestamp 1644511149
transform 1 0 6900 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0579_
timestamp 1644511149
transform -1 0 8096 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0580_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 8280 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0581_
timestamp 1644511149
transform 1 0 8924 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0582_
timestamp 1644511149
transform -1 0 13524 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__or4_2  _0583_
timestamp 1644511149
transform 1 0 19228 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _0584_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 19228 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _0585_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19228 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0586_
timestamp 1644511149
transform -1 0 18860 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0587_
timestamp 1644511149
transform 1 0 16100 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or4_2  _0588_
timestamp 1644511149
transform 1 0 16744 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0589_
timestamp 1644511149
transform -1 0 18032 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0590_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 20700 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0591_
timestamp 1644511149
transform -1 0 20976 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0592_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 18584 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0593_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 18768 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0594_
timestamp 1644511149
transform 1 0 10304 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _0595_
timestamp 1644511149
transform 1 0 13340 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0596_
timestamp 1644511149
transform 1 0 13524 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0597_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11500 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0598_
timestamp 1644511149
transform 1 0 12420 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0599_
timestamp 1644511149
transform -1 0 13340 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0600_
timestamp 1644511149
transform 1 0 11684 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0601_
timestamp 1644511149
transform -1 0 13340 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _0602_
timestamp 1644511149
transform 1 0 10764 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0603_
timestamp 1644511149
transform 1 0 12144 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _0604_
timestamp 1644511149
transform -1 0 9568 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0605_
timestamp 1644511149
transform 1 0 6808 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0606_
timestamp 1644511149
transform 1 0 12788 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0607_
timestamp 1644511149
transform 1 0 14076 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0608_
timestamp 1644511149
transform 1 0 13156 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _0609_
timestamp 1644511149
transform 1 0 13432 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0610_
timestamp 1644511149
transform -1 0 16100 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0611_
timestamp 1644511149
transform 1 0 11132 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _0612_
timestamp 1644511149
transform 1 0 12512 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0613_
timestamp 1644511149
transform 1 0 11868 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0614_
timestamp 1644511149
transform 1 0 13064 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0615_
timestamp 1644511149
transform 1 0 7728 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o41a_1  _0616_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 12052 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0617_
timestamp 1644511149
transform 1 0 12236 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _0618_
timestamp 1644511149
transform 1 0 11684 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0619_
timestamp 1644511149
transform 1 0 9752 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0620_
timestamp 1644511149
transform -1 0 17204 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0621_
timestamp 1644511149
transform 1 0 13340 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _0622_
timestamp 1644511149
transform -1 0 11960 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _0623_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 10580 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0624_
timestamp 1644511149
transform 1 0 19596 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0625_
timestamp 1644511149
transform -1 0 13524 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0626_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 9660 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _0627_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11500 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0628_
timestamp 1644511149
transform -1 0 14720 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0629_
timestamp 1644511149
transform 1 0 14076 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0630_
timestamp 1644511149
transform -1 0 14536 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0631_
timestamp 1644511149
transform 1 0 11500 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0632_
timestamp 1644511149
transform -1 0 12420 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__o31ai_1  _0633_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 10028 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0634_
timestamp 1644511149
transform 1 0 8556 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0635_
timestamp 1644511149
transform 1 0 13616 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _0636_
timestamp 1644511149
transform -1 0 14260 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0637_
timestamp 1644511149
transform 1 0 10764 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _0638_
timestamp 1644511149
transform 1 0 10672 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0639_
timestamp 1644511149
transform 1 0 9936 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _0640_
timestamp 1644511149
transform 1 0 12236 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__or4_2  _0641_
timestamp 1644511149
transform 1 0 14996 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0642_
timestamp 1644511149
transform 1 0 14444 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0643_
timestamp 1644511149
transform -1 0 14996 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _0644_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 12696 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _0645_
timestamp 1644511149
transform 1 0 12512 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _0646_
timestamp 1644511149
transform 1 0 9016 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0647_
timestamp 1644511149
transform -1 0 16836 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0648_
timestamp 1644511149
transform 1 0 16652 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0649_
timestamp 1644511149
transform 1 0 16100 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0650_
timestamp 1644511149
transform 1 0 17388 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0651_
timestamp 1644511149
transform -1 0 13064 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0652_
timestamp 1644511149
transform 1 0 9476 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _0653_
timestamp 1644511149
transform 1 0 9568 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0654_
timestamp 1644511149
transform -1 0 9936 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0655_
timestamp 1644511149
transform -1 0 12604 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _0656_
timestamp 1644511149
transform 1 0 10120 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_2  _0657_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 17204 0 1 9792
box -38 -48 1234 592
use sky130_fd_sc_hd__or3_1  _0658_
timestamp 1644511149
transform 1 0 10212 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0659_
timestamp 1644511149
transform -1 0 12788 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__a211o_1  _0660_
timestamp 1644511149
transform 1 0 10672 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0661_
timestamp 1644511149
transform -1 0 13800 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0662_
timestamp 1644511149
transform -1 0 11040 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0663_
timestamp 1644511149
transform 1 0 14076 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__o21ai_1  _0664_
timestamp 1644511149
transform 1 0 13616 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _0665_
timestamp 1644511149
transform 1 0 15180 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__or4_2  _0666_
timestamp 1644511149
transform -1 0 15272 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _0667_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 14996 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0668_
timestamp 1644511149
transform 1 0 13248 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0669_
timestamp 1644511149
transform 1 0 14168 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _0670_
timestamp 1644511149
transform -1 0 12788 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0671_
timestamp 1644511149
transform 1 0 10948 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _0672_
timestamp 1644511149
transform 1 0 11868 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0673_
timestamp 1644511149
transform -1 0 20240 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0674_
timestamp 1644511149
transform 1 0 11684 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0675_
timestamp 1644511149
transform 1 0 11408 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0676_
timestamp 1644511149
transform -1 0 12788 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _0677_
timestamp 1644511149
transform -1 0 15364 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _0678_
timestamp 1644511149
transform -1 0 12144 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _0679_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 12236 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _0680_
timestamp 1644511149
transform 1 0 12052 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0681_
timestamp 1644511149
transform -1 0 11868 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _0682_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 15640 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0683_
timestamp 1644511149
transform -1 0 13524 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _0684_
timestamp 1644511149
transform 1 0 12052 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0685_
timestamp 1644511149
transform 1 0 10856 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _0686_
timestamp 1644511149
transform 1 0 12880 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _0687_
timestamp 1644511149
transform 1 0 12972 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0688_
timestamp 1644511149
transform -1 0 13800 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0689_
timestamp 1644511149
transform 1 0 6992 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0690_
timestamp 1644511149
transform 1 0 6900 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0691_
timestamp 1644511149
transform 1 0 7912 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0692_
timestamp 1644511149
transform 1 0 9384 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0693_
timestamp 1644511149
transform 1 0 9292 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0694_
timestamp 1644511149
transform 1 0 9384 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0695_
timestamp 1644511149
transform 1 0 7820 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0696_
timestamp 1644511149
transform 1 0 7176 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0697_
timestamp 1644511149
transform -1 0 8096 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0698_
timestamp 1644511149
transform 1 0 7820 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0699_
timestamp 1644511149
transform -1 0 7636 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0700_
timestamp 1644511149
transform -1 0 6992 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0701_
timestamp 1644511149
transform 1 0 8924 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0702_
timestamp 1644511149
transform 1 0 8648 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0703_
timestamp 1644511149
transform 1 0 9292 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0704_
timestamp 1644511149
transform -1 0 13800 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _0705_
timestamp 1644511149
transform 1 0 7452 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0706_
timestamp 1644511149
transform 1 0 6716 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0707_
timestamp 1644511149
transform 1 0 6808 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0708_
timestamp 1644511149
transform 1 0 6992 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0709_
timestamp 1644511149
transform -1 0 6808 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0710_
timestamp 1644511149
transform -1 0 6072 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0711_
timestamp 1644511149
transform 1 0 7268 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0712_
timestamp 1644511149
transform 1 0 6624 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0713_
timestamp 1644511149
transform 1 0 8280 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0714_
timestamp 1644511149
transform 1 0 7268 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0715_
timestamp 1644511149
transform -1 0 6072 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0716_
timestamp 1644511149
transform -1 0 5428 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0717_
timestamp 1644511149
transform -1 0 6900 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0718_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 8924 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0719_
timestamp 1644511149
transform 1 0 7728 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _0720_
timestamp 1644511149
transform 1 0 7360 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0721_
timestamp 1644511149
transform 1 0 10764 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0722_
timestamp 1644511149
transform -1 0 11316 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0723_
timestamp 1644511149
transform -1 0 9016 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0724_
timestamp 1644511149
transform 1 0 9752 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0725_
timestamp 1644511149
transform -1 0 10396 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0726_
timestamp 1644511149
transform 1 0 9660 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__o31ai_1  _0727_
timestamp 1644511149
transform 1 0 9476 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0728_
timestamp 1644511149
transform -1 0 22080 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0729_
timestamp 1644511149
transform 1 0 21160 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _0730_
timestamp 1644511149
transform -1 0 10948 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0731_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 8648 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _0732_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 8280 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0733_
timestamp 1644511149
transform -1 0 19596 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _0734_
timestamp 1644511149
transform 1 0 7084 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0735_
timestamp 1644511149
transform -1 0 9384 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0736_
timestamp 1644511149
transform -1 0 8924 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0737_
timestamp 1644511149
transform -1 0 9200 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0738_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 8648 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0739_
timestamp 1644511149
transform 1 0 23276 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a2111oi_1  _0740_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 8004 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _0741_
timestamp 1644511149
transform -1 0 10304 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_1  _0742_
timestamp 1644511149
transform 1 0 8924 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _0743_
timestamp 1644511149
transform -1 0 9660 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0744_
timestamp 1644511149
transform 1 0 7912 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0745_
timestamp 1644511149
transform -1 0 9200 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0746_
timestamp 1644511149
transform -1 0 7728 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0747_
timestamp 1644511149
transform -1 0 7636 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0748_
timestamp 1644511149
transform 1 0 6900 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0749_
timestamp 1644511149
transform -1 0 7636 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0750_
timestamp 1644511149
transform -1 0 7268 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a2111oi_1  _0751_
timestamp 1644511149
transform 1 0 6256 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _0752_
timestamp 1644511149
transform 1 0 6532 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0753_
timestamp 1644511149
transform 1 0 7544 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0754_
timestamp 1644511149
transform 1 0 5520 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0755_
timestamp 1644511149
transform -1 0 5428 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a311o_1  _0756_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6532 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _0757_
timestamp 1644511149
transform 1 0 5612 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _0758_
timestamp 1644511149
transform -1 0 20884 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0759_
timestamp 1644511149
transform 1 0 19228 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _0760_
timestamp 1644511149
transform -1 0 18492 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0761_
timestamp 1644511149
transform -1 0 20332 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0762_
timestamp 1644511149
transform 1 0 19044 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0763_
timestamp 1644511149
transform -1 0 21528 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0764_
timestamp 1644511149
transform -1 0 22632 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0765_
timestamp 1644511149
transform 1 0 17848 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__or2b_1  _0766_
timestamp 1644511149
transform -1 0 18308 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0767_
timestamp 1644511149
transform -1 0 19872 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0768_
timestamp 1644511149
transform 1 0 19228 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__nand3b_2  _0769_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16652 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__or4_2  _0770_
timestamp 1644511149
transform -1 0 16376 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0771_
timestamp 1644511149
transform 1 0 15364 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__nor4_2  _0772_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 17940 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__nor4_2  _0773_
timestamp 1644511149
transform -1 0 17572 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _0774_
timestamp 1644511149
transform 1 0 14904 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__and4bb_1  _0775_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 19596 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _0776_
timestamp 1644511149
transform -1 0 12420 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0777_
timestamp 1644511149
transform 1 0 19780 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0778_
timestamp 1644511149
transform -1 0 11960 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0779_
timestamp 1644511149
transform 1 0 12604 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _0780_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14076 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0781_
timestamp 1644511149
transform -1 0 22724 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0782_
timestamp 1644511149
transform 1 0 21252 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0783_
timestamp 1644511149
transform -1 0 20792 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0784_
timestamp 1644511149
transform 1 0 13800 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _0785_
timestamp 1644511149
transform 1 0 12880 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0786_
timestamp 1644511149
transform 1 0 16652 0 -1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0787_
timestamp 1644511149
transform -1 0 16376 0 -1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _0788_
timestamp 1644511149
transform 1 0 15824 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _0789_
timestamp 1644511149
transform 1 0 13800 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0790_
timestamp 1644511149
transform -1 0 20700 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0791_
timestamp 1644511149
transform 1 0 14076 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _0792_
timestamp 1644511149
transform 1 0 12236 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0793_
timestamp 1644511149
transform 1 0 15088 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _0794_
timestamp 1644511149
transform -1 0 15640 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0795_
timestamp 1644511149
transform 1 0 21068 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0796_
timestamp 1644511149
transform -1 0 21988 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _0797_
timestamp 1644511149
transform 1 0 13156 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0798_
timestamp 1644511149
transform 1 0 15732 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _0799_
timestamp 1644511149
transform 1 0 14628 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0800_
timestamp 1644511149
transform -1 0 22080 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0801_
timestamp 1644511149
transform 1 0 14076 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _0802_
timestamp 1644511149
transform 1 0 13248 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0803_
timestamp 1644511149
transform 1 0 15916 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _0804_
timestamp 1644511149
transform -1 0 16008 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0805_
timestamp 1644511149
transform 1 0 22172 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0806_
timestamp 1644511149
transform -1 0 21252 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _0807_
timestamp 1644511149
transform -1 0 22540 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _0808_
timestamp 1644511149
transform 1 0 13248 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0809_
timestamp 1644511149
transform 1 0 16652 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _0810_
timestamp 1644511149
transform -1 0 16284 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0811_
timestamp 1644511149
transform -1 0 22264 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0812_
timestamp 1644511149
transform -1 0 22448 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _0813_
timestamp 1644511149
transform 1 0 13340 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0814_
timestamp 1644511149
transform -1 0 13800 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _0815_
timestamp 1644511149
transform -1 0 15456 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0816_
timestamp 1644511149
transform 1 0 21712 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0817_
timestamp 1644511149
transform -1 0 22540 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _0818_
timestamp 1644511149
transform 1 0 12604 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0819_
timestamp 1644511149
transform 1 0 12512 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _0820_
timestamp 1644511149
transform -1 0 14628 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0821_
timestamp 1644511149
transform -1 0 21436 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0822_
timestamp 1644511149
transform 1 0 20608 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0823_
timestamp 1644511149
transform 1 0 6348 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _0824_
timestamp 1644511149
transform 1 0 7636 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0825_
timestamp 1644511149
transform -1 0 7820 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0826_
timestamp 1644511149
transform -1 0 8096 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0827_
timestamp 1644511149
transform 1 0 7360 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0828_
timestamp 1644511149
transform 1 0 8004 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _0829_
timestamp 1644511149
transform 1 0 7728 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _0830_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6440 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _0831_
timestamp 1644511149
transform 1 0 5796 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0832_
timestamp 1644511149
transform -1 0 8280 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _0833_
timestamp 1644511149
transform 1 0 6348 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__o31ai_1  _0834_
timestamp 1644511149
transform -1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0835_
timestamp 1644511149
transform -1 0 7176 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0836_
timestamp 1644511149
transform -1 0 15180 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0837_
timestamp 1644511149
transform 1 0 15548 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0838_
timestamp 1644511149
transform 1 0 14536 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0839_
timestamp 1644511149
transform 1 0 13248 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0840_
timestamp 1644511149
transform -1 0 13984 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0841_
timestamp 1644511149
transform -1 0 15364 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _0842_
timestamp 1644511149
transform -1 0 16928 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0843_
timestamp 1644511149
transform -1 0 17572 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0844_
timestamp 1644511149
transform -1 0 15916 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0845_
timestamp 1644511149
transform 1 0 16192 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0846_
timestamp 1644511149
transform 1 0 15548 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0847_
timestamp 1644511149
transform -1 0 18032 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0848_
timestamp 1644511149
transform 1 0 16192 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0849_
timestamp 1644511149
transform 1 0 15916 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0850_
timestamp 1644511149
transform -1 0 16928 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0851_
timestamp 1644511149
transform 1 0 14904 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0852_
timestamp 1644511149
transform 1 0 14260 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0853_
timestamp 1644511149
transform 1 0 14720 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0854_
timestamp 1644511149
transform -1 0 15548 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0855_
timestamp 1644511149
transform 1 0 15732 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0856_
timestamp 1644511149
transform 1 0 16652 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0857_
timestamp 1644511149
transform 1 0 19596 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _0858_
timestamp 1644511149
transform -1 0 15088 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0859_
timestamp 1644511149
transform 1 0 20700 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _0860_
timestamp 1644511149
transform 1 0 14536 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0861_
timestamp 1644511149
transform 1 0 14076 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _0862_
timestamp 1644511149
transform 1 0 16008 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _0863_
timestamp 1644511149
transform -1 0 16652 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0864_
timestamp 1644511149
transform 1 0 14076 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0865_
timestamp 1644511149
transform -1 0 18492 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0866_
timestamp 1644511149
transform -1 0 16192 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0867_
timestamp 1644511149
transform -1 0 17112 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0868_
timestamp 1644511149
transform 1 0 17296 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0869_
timestamp 1644511149
transform -1 0 15364 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0870_
timestamp 1644511149
transform 1 0 15088 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0871_
timestamp 1644511149
transform 1 0 17940 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _0872_
timestamp 1644511149
transform 1 0 16652 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0873_
timestamp 1644511149
transform -1 0 17664 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _0874_
timestamp 1644511149
transform 1 0 17388 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a2111o_1  _0875_
timestamp 1644511149
transform 1 0 17940 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _0876_
timestamp 1644511149
transform 1 0 17204 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__or4_2  _0877_
timestamp 1644511149
transform -1 0 19412 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0878_
timestamp 1644511149
transform -1 0 18400 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0879_
timestamp 1644511149
transform 1 0 17204 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0880_
timestamp 1644511149
transform -1 0 16928 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0881_
timestamp 1644511149
transform 1 0 17664 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _0882_
timestamp 1644511149
transform -1 0 17480 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_1  _0883_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 15640 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _0884_
timestamp 1644511149
transform 1 0 16100 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0885_
timestamp 1644511149
transform -1 0 17020 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _0886_
timestamp 1644511149
transform 1 0 18952 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__o31ai_1  _0887_
timestamp 1644511149
transform 1 0 19228 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0888_
timestamp 1644511149
transform 1 0 18584 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a221oi_1  _0889_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 19872 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0890_
timestamp 1644511149
transform 1 0 23276 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _0891_
timestamp 1644511149
transform 1 0 19964 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0892_
timestamp 1644511149
transform 1 0 21804 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a211oi_1  _0893_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 23092 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _0894_
timestamp 1644511149
transform 1 0 21344 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0895_
timestamp 1644511149
transform 1 0 23092 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0896_
timestamp 1644511149
transform 1 0 20608 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0897_
timestamp 1644511149
transform -1 0 5888 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0898_
timestamp 1644511149
transform 1 0 5428 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0899_
timestamp 1644511149
transform 1 0 24380 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _0900_
timestamp 1644511149
transform -1 0 24012 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0901_
timestamp 1644511149
transform -1 0 24104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0902_
timestamp 1644511149
transform -1 0 16744 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0903_
timestamp 1644511149
transform 1 0 16652 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _0904_
timestamp 1644511149
transform 1 0 16008 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__nor4_1  _0905_
timestamp 1644511149
transform -1 0 16376 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0906_
timestamp 1644511149
transform -1 0 16008 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0907_
timestamp 1644511149
transform 1 0 16744 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0908_
timestamp 1644511149
transform -1 0 17940 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0909_
timestamp 1644511149
transform -1 0 14628 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0910_
timestamp 1644511149
transform -1 0 21344 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _0911_
timestamp 1644511149
transform 1 0 14168 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0912_
timestamp 1644511149
transform 1 0 14812 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0913_
timestamp 1644511149
transform 1 0 15088 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0914_
timestamp 1644511149
transform 1 0 15916 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _0915_
timestamp 1644511149
transform -1 0 16652 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0916_
timestamp 1644511149
transform 1 0 17388 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0917_
timestamp 1644511149
transform -1 0 17848 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0918_
timestamp 1644511149
transform -1 0 13800 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0919_
timestamp 1644511149
transform 1 0 14076 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0920_
timestamp 1644511149
transform -1 0 14352 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0921_
timestamp 1644511149
transform 1 0 13432 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0922_
timestamp 1644511149
transform -1 0 15548 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0923_
timestamp 1644511149
transform -1 0 21528 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _0924_
timestamp 1644511149
transform 1 0 14996 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__and4b_1  _0925_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17664 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0926_
timestamp 1644511149
transform 1 0 18400 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or3_2  _0927_
timestamp 1644511149
transform 1 0 19228 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0928_
timestamp 1644511149
transform 1 0 19228 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _0929_
timestamp 1644511149
transform -1 0 18860 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0930_
timestamp 1644511149
transform -1 0 18400 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0931_
timestamp 1644511149
transform -1 0 19688 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0932_
timestamp 1644511149
transform 1 0 19412 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0933_
timestamp 1644511149
transform 1 0 19872 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0934_
timestamp 1644511149
transform 1 0 19964 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0935_
timestamp 1644511149
transform -1 0 21160 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0936_
timestamp 1644511149
transform 1 0 19964 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0937_
timestamp 1644511149
transform 1 0 19320 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0938_
timestamp 1644511149
transform -1 0 21160 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0939_
timestamp 1644511149
transform -1 0 18952 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0940_
timestamp 1644511149
transform -1 0 19596 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0941_
timestamp 1644511149
transform 1 0 18216 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0942_
timestamp 1644511149
transform 1 0 19228 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0943_
timestamp 1644511149
transform 1 0 18492 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0944_
timestamp 1644511149
transform 1 0 18676 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0945_
timestamp 1644511149
transform 1 0 20240 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0946_
timestamp 1644511149
transform 1 0 20056 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0947_
timestamp 1644511149
transform 1 0 21252 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0948_
timestamp 1644511149
transform 1 0 12144 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _0949_
timestamp 1644511149
transform 1 0 14536 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0950_
timestamp 1644511149
transform 1 0 12236 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0951_
timestamp 1644511149
transform -1 0 13064 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0952_
timestamp 1644511149
transform 1 0 13524 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0953_
timestamp 1644511149
transform 1 0 12512 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0954_
timestamp 1644511149
transform 1 0 13248 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0955_
timestamp 1644511149
transform 1 0 17572 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__or2b_1  _0956_
timestamp 1644511149
transform 1 0 17020 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _0957_
timestamp 1644511149
transform -1 0 17940 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__nor4_1  _0958_
timestamp 1644511149
transform -1 0 18216 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0959_
timestamp 1644511149
transform 1 0 20516 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0960_
timestamp 1644511149
transform 1 0 22908 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0961_
timestamp 1644511149
transform -1 0 23000 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0962_
timestamp 1644511149
transform 1 0 22356 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0963_
timestamp 1644511149
transform -1 0 23552 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _0964_
timestamp 1644511149
transform -1 0 21344 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0965_
timestamp 1644511149
transform 1 0 20240 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0966_
timestamp 1644511149
transform -1 0 19872 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0967_
timestamp 1644511149
transform 1 0 20056 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0968_
timestamp 1644511149
transform -1 0 23276 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0969_
timestamp 1644511149
transform -1 0 22632 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0970_
timestamp 1644511149
transform 1 0 22908 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0971_
timestamp 1644511149
transform 1 0 22264 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _0972_
timestamp 1644511149
transform -1 0 23552 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0973_
timestamp 1644511149
transform 1 0 23460 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0974_
timestamp 1644511149
transform -1 0 23920 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0975_
timestamp 1644511149
transform -1 0 24012 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0976_
timestamp 1644511149
transform -1 0 23920 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0977_
timestamp 1644511149
transform -1 0 23828 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0978_
timestamp 1644511149
transform -1 0 23736 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0979_
timestamp 1644511149
transform 1 0 24380 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0980_
timestamp 1644511149
transform -1 0 23736 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0981_
timestamp 1644511149
transform 1 0 11500 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0982_
timestamp 1644511149
transform 1 0 10764 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0983_
timestamp 1644511149
transform -1 0 11684 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0984_
timestamp 1644511149
transform 1 0 11776 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0985_
timestamp 1644511149
transform 1 0 10764 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0986_
timestamp 1644511149
transform -1 0 11224 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0987_
timestamp 1644511149
transform -1 0 11408 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0988_
timestamp 1644511149
transform 1 0 10396 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0989_
timestamp 1644511149
transform 1 0 10120 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0990_
timestamp 1644511149
transform 1 0 11500 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0991_
timestamp 1644511149
transform 1 0 10948 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0992_
timestamp 1644511149
transform 1 0 10396 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0993_
timestamp 1644511149
transform 1 0 10396 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0994_
timestamp 1644511149
transform -1 0 11224 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0995_
timestamp 1644511149
transform 1 0 9108 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0996_
timestamp 1644511149
transform -1 0 9384 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0997_
timestamp 1644511149
transform -1 0 8740 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0998_
timestamp 1644511149
transform 1 0 10304 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0999_
timestamp 1644511149
transform 1 0 10396 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1000_
timestamp 1644511149
transform -1 0 11684 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1001_
timestamp 1644511149
transform 1 0 9200 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1002_
timestamp 1644511149
transform 1 0 8648 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1003_
timestamp 1644511149
transform -1 0 9752 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1004_
timestamp 1644511149
transform 1 0 11500 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1005_
timestamp 1644511149
transform 1 0 11040 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1006_
timestamp 1644511149
transform -1 0 12604 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1007_
timestamp 1644511149
transform -1 0 21804 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1008_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 19228 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__or4b_2  _1009_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 18216 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1010_
timestamp 1644511149
transform 1 0 21804 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1011_
timestamp 1644511149
transform -1 0 25300 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1012_
timestamp 1644511149
transform 1 0 24748 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1013_
timestamp 1644511149
transform -1 0 25668 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1014_
timestamp 1644511149
transform 1 0 19872 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1015_
timestamp 1644511149
transform -1 0 20148 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1016_
timestamp 1644511149
transform -1 0 19596 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1017_
timestamp 1644511149
transform 1 0 22172 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1018_
timestamp 1644511149
transform 1 0 21528 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1019_
timestamp 1644511149
transform 1 0 23000 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1020_
timestamp 1644511149
transform 1 0 20056 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1021_
timestamp 1644511149
transform 1 0 20332 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1022_
timestamp 1644511149
transform -1 0 19044 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1023_
timestamp 1644511149
transform 1 0 24380 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1024_
timestamp 1644511149
transform 1 0 24380 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1025_
timestamp 1644511149
transform 1 0 25852 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1026_
timestamp 1644511149
transform 1 0 23644 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1027_
timestamp 1644511149
transform 1 0 23460 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1028_
timestamp 1644511149
transform -1 0 24104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1029_
timestamp 1644511149
transform 1 0 20424 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1030_
timestamp 1644511149
transform 1 0 20332 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1031_
timestamp 1644511149
transform 1 0 21068 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1032_
timestamp 1644511149
transform 1 0 22172 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1033_
timestamp 1644511149
transform 1 0 21804 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1034_
timestamp 1644511149
transform 1 0 23368 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1035_
timestamp 1644511149
transform 1 0 19964 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1036_
timestamp 1644511149
transform -1 0 25852 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1037_
timestamp 1644511149
transform 1 0 24380 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1038_
timestamp 1644511149
transform 1 0 22632 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a211oi_1  _1039_
timestamp 1644511149
transform -1 0 23460 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a211oi_1  _1040_
timestamp 1644511149
transform 1 0 21804 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a311oi_1  _1041_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20792 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1042_
timestamp 1644511149
transform -1 0 22264 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1043_
timestamp 1644511149
transform -1 0 22448 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _1044_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 20608 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1045_
timestamp 1644511149
transform 1 0 20884 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1046_
timestamp 1644511149
transform 1 0 20056 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1047_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 9476 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1048_
timestamp 1644511149
transform -1 0 18032 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1049_
timestamp 1644511149
transform 1 0 8924 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1050_
timestamp 1644511149
transform 1 0 8372 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1051_
timestamp 1644511149
transform 1 0 9476 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1052_
timestamp 1644511149
transform 1 0 12144 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1053_
timestamp 1644511149
transform 1 0 7912 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1054_
timestamp 1644511149
transform 1 0 8372 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1055_
timestamp 1644511149
transform -1 0 15456 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1056_
timestamp 1644511149
transform 1 0 12144 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1057_
timestamp 1644511149
transform 1 0 11684 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1058_
timestamp 1644511149
transform -1 0 14812 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1059_
timestamp 1644511149
transform 1 0 9292 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1060_
timestamp 1644511149
transform 1 0 7636 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1061_
timestamp 1644511149
transform 1 0 6808 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1062_
timestamp 1644511149
transform 1 0 9016 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1063_
timestamp 1644511149
transform 1 0 6624 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1064_
timestamp 1644511149
transform 1 0 5980 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1065_
timestamp 1644511149
transform -1 0 8648 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1066_
timestamp 1644511149
transform 1 0 5612 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1067_
timestamp 1644511149
transform 1 0 11500 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1068_
timestamp 1644511149
transform -1 0 12052 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1069_
timestamp 1644511149
transform 1 0 9108 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1070_
timestamp 1644511149
transform 1 0 7820 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1071_
timestamp 1644511149
transform 1 0 9476 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1072_
timestamp 1644511149
transform 1 0 6532 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1073_
timestamp 1644511149
transform 1 0 4600 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1074_
timestamp 1644511149
transform 1 0 4416 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1075_
timestamp 1644511149
transform -1 0 5980 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1076_
timestamp 1644511149
transform -1 0 7912 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1077_
timestamp 1644511149
transform -1 0 6072 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1078_
timestamp 1644511149
transform 1 0 22080 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1079_
timestamp 1644511149
transform -1 0 8188 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1080_
timestamp 1644511149
transform 1 0 22632 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1081_
timestamp 1644511149
transform 1 0 23736 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1082_
timestamp 1644511149
transform 1 0 24380 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1083_
timestamp 1644511149
transform 1 0 20700 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1084_
timestamp 1644511149
transform 1 0 4600 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1085_
timestamp 1644511149
transform -1 0 6716 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1086_
timestamp 1644511149
transform 1 0 4600 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1087_
timestamp 1644511149
transform 1 0 5980 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1088_
timestamp 1644511149
transform 1 0 14076 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1089_
timestamp 1644511149
transform 1 0 16652 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1090_
timestamp 1644511149
transform -1 0 18124 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1091_
timestamp 1644511149
transform 1 0 16652 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1092_
timestamp 1644511149
transform 1 0 14352 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1093_
timestamp 1644511149
transform -1 0 15732 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1094_
timestamp 1644511149
transform 1 0 14076 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1095_
timestamp 1644511149
transform 1 0 15732 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1096_
timestamp 1644511149
transform 1 0 14904 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1097_
timestamp 1644511149
transform 1 0 17480 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1098_
timestamp 1644511149
transform 1 0 17756 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1099_
timestamp 1644511149
transform 1 0 16652 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1100_
timestamp 1644511149
transform 1 0 16192 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1101_
timestamp 1644511149
transform 1 0 18952 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1102_
timestamp 1644511149
transform -1 0 24288 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1103_
timestamp 1644511149
transform 1 0 20056 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1104_
timestamp 1644511149
transform 1 0 5152 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1105_
timestamp 1644511149
transform 1 0 25208 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1106_
timestamp 1644511149
transform 1 0 25208 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1107_
timestamp 1644511149
transform 1 0 23460 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1108_
timestamp 1644511149
transform 1 0 22632 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1109_
timestamp 1644511149
transform -1 0 27048 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1110_
timestamp 1644511149
transform 1 0 25760 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1111_
timestamp 1644511149
transform 1 0 23460 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1112_
timestamp 1644511149
transform 1 0 21344 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1113_
timestamp 1644511149
transform -1 0 23276 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1114_
timestamp 1644511149
transform 1 0 23736 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1115_
timestamp 1644511149
transform -1 0 18952 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1116_
timestamp 1644511149
transform 1 0 14076 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1117_
timestamp 1644511149
transform -1 0 13800 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1118_
timestamp 1644511149
transform -1 0 18124 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1119_
timestamp 1644511149
transform -1 0 18860 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1120_
timestamp 1644511149
transform 1 0 11316 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1121_
timestamp 1644511149
transform 1 0 14352 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1122_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14076 0 1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1123_
timestamp 1644511149
transform 1 0 18216 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1124_
timestamp 1644511149
transform -1 0 23276 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1125_
timestamp 1644511149
transform -1 0 22448 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1126_
timestamp 1644511149
transform 1 0 17480 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1127_
timestamp 1644511149
transform 1 0 18308 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1128_
timestamp 1644511149
transform -1 0 21528 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1129_
timestamp 1644511149
transform 1 0 12880 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1130_
timestamp 1644511149
transform 1 0 12328 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1131_
timestamp 1644511149
transform 1 0 17480 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1132_
timestamp 1644511149
transform 1 0 18032 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1133_
timestamp 1644511149
transform 1 0 19596 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1134_
timestamp 1644511149
transform -1 0 20700 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1135_
timestamp 1644511149
transform 1 0 22356 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1136_
timestamp 1644511149
transform 1 0 23736 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1137_
timestamp 1644511149
transform 1 0 24380 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1138_
timestamp 1644511149
transform 1 0 23920 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1139_
timestamp 1644511149
transform 1 0 24380 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1140_
timestamp 1644511149
transform 1 0 23920 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1141_
timestamp 1644511149
transform -1 0 12144 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1142_
timestamp 1644511149
transform 1 0 11868 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1143_
timestamp 1644511149
transform 1 0 10948 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1144_
timestamp 1644511149
transform 1 0 11500 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1145_
timestamp 1644511149
transform 1 0 8924 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1146_
timestamp 1644511149
transform 1 0 11500 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1147_
timestamp 1644511149
transform 1 0 9292 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1148_
timestamp 1644511149
transform -1 0 13156 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1149_
timestamp 1644511149
transform 1 0 25484 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1150_
timestamp 1644511149
transform 1 0 19780 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1151_
timestamp 1644511149
transform 1 0 22356 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1152_
timestamp 1644511149
transform 1 0 19596 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1153_
timestamp 1644511149
transform 1 0 25392 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1154_
timestamp 1644511149
transform -1 0 25852 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1155_
timestamp 1644511149
transform 1 0 20056 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1156_
timestamp 1644511149
transform -1 0 23276 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1157_
timestamp 1644511149
transform 1 0 26036 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1158_
timestamp 1644511149
transform 1 0 22632 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1159_
timestamp 1644511149
transform -1 0 23092 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1160_
timestamp 1644511149
transform 1 0 19964 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1161_
timestamp 1644511149
transform 1 0 19688 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _1162__33 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 28152 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1163__34
timestamp 1644511149
transform 1 0 28152 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1164__35
timestamp 1644511149
transform -1 0 19688 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1165__36
timestamp 1644511149
transform -1 0 1656 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1166__37
timestamp 1644511149
transform -1 0 1656 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1167__38
timestamp 1644511149
transform 1 0 28152 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1168__39
timestamp 1644511149
transform -1 0 1656 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1169__40
timestamp 1644511149
transform -1 0 1656 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1170__41
timestamp 1644511149
transform 1 0 28152 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1171__42
timestamp 1644511149
transform -1 0 1656 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1172__43
timestamp 1644511149
transform 1 0 28152 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1173__44
timestamp 1644511149
transform -1 0 1656 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1174__45
timestamp 1644511149
transform -1 0 26128 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1175__46
timestamp 1644511149
transform -1 0 27232 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1176__47
timestamp 1644511149
transform 1 0 28152 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1177__48
timestamp 1644511149
transform 1 0 28152 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1178__49
timestamp 1644511149
transform 1 0 28152 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1179__50
timestamp 1644511149
transform -1 0 4232 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1180__51
timestamp 1644511149
transform -1 0 1656 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1181__52
timestamp 1644511149
transform -1 0 22080 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1182__53
timestamp 1644511149
transform -1 0 12604 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1183__54
timestamp 1644511149
transform 1 0 27600 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1184__55
timestamp 1644511149
transform -1 0 6808 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1185__56
timestamp 1644511149
transform -1 0 4048 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clock pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 15824 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_0_0_clock
timestamp 1644511149
transform -1 0 10212 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_1_0_clock
timestamp 1644511149
transform 1 0 11500 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_2_0_clock
timestamp 1644511149
transform -1 0 21988 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_3_0_clock
timestamp 1644511149
transform 1 0 21988 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_4_0_clock
timestamp 1644511149
transform 1 0 9660 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_5_0_clock
timestamp 1644511149
transform -1 0 10488 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_6_0_clock
timestamp 1644511149
transform -1 0 21804 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_7_0_clock
timestamp 1644511149
transform -1 0 19688 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_0_0_clock
timestamp 1644511149
transform -1 0 9476 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_1_0_clock
timestamp 1644511149
transform 1 0 11500 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_2_0_clock
timestamp 1644511149
transform -1 0 9292 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_3_0_clock
timestamp 1644511149
transform 1 0 11960 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_4_0_clock
timestamp 1644511149
transform -1 0 19872 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_5_0_clock
timestamp 1644511149
transform 1 0 23276 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_6_0_clock
timestamp 1644511149
transform -1 0 19504 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_7_0_clock
timestamp 1644511149
transform 1 0 23460 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_8_0_clock
timestamp 1644511149
transform -1 0 8832 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_9_0_clock
timestamp 1644511149
transform 1 0 11592 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_10_0_clock
timestamp 1644511149
transform -1 0 9108 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_11_0_clock
timestamp 1644511149
transform 1 0 13156 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_12_0_clock
timestamp 1644511149
transform -1 0 18952 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_13_0_clock
timestamp 1644511149
transform 1 0 24104 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_14_0_clock
timestamp 1644511149
transform -1 0 17572 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_15_0_clock
timestamp 1644511149
transform 1 0 20608 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input1
timestamp 1644511149
transform 1 0 1380 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  input2 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 1564 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input3
timestamp 1644511149
transform 1 0 10396 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input4
timestamp 1644511149
transform -1 0 28428 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input5
timestamp 1644511149
transform 1 0 19228 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input6
timestamp 1644511149
transform -1 0 28152 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input7
timestamp 1644511149
transform 1 0 1564 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1644511149
transform 1 0 28152 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1644511149
transform 1 0 20700 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input10
timestamp 1644511149
transform 1 0 1380 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input11
timestamp 1644511149
transform -1 0 28428 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input12
timestamp 1644511149
transform 1 0 1564 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input13
timestamp 1644511149
transform 1 0 5244 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input14
timestamp 1644511149
transform -1 0 28428 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input15
timestamp 1644511149
transform 1 0 16836 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input16
timestamp 1644511149
transform 1 0 24564 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input17
timestamp 1644511149
transform 1 0 22632 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input18
timestamp 1644511149
transform 1 0 2668 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input19
timestamp 1644511149
transform 1 0 1564 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input20
timestamp 1644511149
transform 1 0 1380 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input21
timestamp 1644511149
transform -1 0 28428 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output22
timestamp 1644511149
transform 1 0 25208 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output23
timestamp 1644511149
transform -1 0 17020 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output24
timestamp 1644511149
transform 1 0 28060 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output25
timestamp 1644511149
transform -1 0 2484 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output26
timestamp 1644511149
transform -1 0 1748 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output27
timestamp 1644511149
transform 1 0 28060 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output28
timestamp 1644511149
transform -1 0 1748 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output29
timestamp 1644511149
transform 1 0 28060 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output30
timestamp 1644511149
transform 1 0 25300 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output31
timestamp 1644511149
transform 1 0 28060 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output32
timestamp 1644511149
transform -1 0 22356 0 1 2176
box -38 -48 406 592
<< labels >>
rlabel metal2 s 9034 29200 9090 30000 6 clock
port 0 nsew signal input
rlabel metal3 s 0 19728 800 19848 6 io_rxd
port 1 nsew signal input
rlabel metal2 s 25134 0 25190 800 6 io_txd
port 2 nsew signal tristate
rlabel metal2 s 16118 29200 16174 30000 6 io_uartInt
port 3 nsew signal tristate
rlabel metal3 s 0 27888 800 28008 6 io_uart_select
port 4 nsew signal input
rlabel metal3 s 29200 10208 30000 10328 6 io_wbs_ack_o
port 5 nsew signal tristate
rlabel metal3 s 0 2048 800 2168 6 io_wbs_data_o[0]
port 6 nsew signal tristate
rlabel metal2 s 19338 29200 19394 30000 6 io_wbs_data_o[10]
port 7 nsew signal tristate
rlabel metal3 s 0 21088 800 21208 6 io_wbs_data_o[11]
port 8 nsew signal tristate
rlabel metal3 s 0 10208 800 10328 6 io_wbs_data_o[12]
port 9 nsew signal tristate
rlabel metal3 s 29200 23128 30000 23248 6 io_wbs_data_o[13]
port 10 nsew signal tristate
rlabel metal3 s 0 23128 800 23248 6 io_wbs_data_o[14]
port 11 nsew signal tristate
rlabel metal3 s 0 17008 800 17128 6 io_wbs_data_o[15]
port 12 nsew signal tristate
rlabel metal3 s 29200 5448 30000 5568 6 io_wbs_data_o[16]
port 13 nsew signal tristate
rlabel metal3 s 0 13608 800 13728 6 io_wbs_data_o[17]
port 14 nsew signal tristate
rlabel metal3 s 29200 14968 30000 15088 6 io_wbs_data_o[18]
port 15 nsew signal tristate
rlabel metal3 s 0 25848 800 25968 6 io_wbs_data_o[19]
port 16 nsew signal tristate
rlabel metal3 s 0 16328 800 16448 6 io_wbs_data_o[1]
port 17 nsew signal tristate
rlabel metal2 s 25778 29200 25834 30000 6 io_wbs_data_o[20]
port 18 nsew signal tristate
rlabel metal2 s 26422 0 26478 800 6 io_wbs_data_o[21]
port 19 nsew signal tristate
rlabel metal3 s 29200 4088 30000 4208 6 io_wbs_data_o[22]
port 20 nsew signal tristate
rlabel metal3 s 29200 16328 30000 16448 6 io_wbs_data_o[23]
port 21 nsew signal tristate
rlabel metal3 s 29200 26528 30000 26648 6 io_wbs_data_o[24]
port 22 nsew signal tristate
rlabel metal2 s 3882 29200 3938 30000 6 io_wbs_data_o[25]
port 23 nsew signal tristate
rlabel metal3 s 0 18368 800 18488 6 io_wbs_data_o[26]
port 24 nsew signal tristate
rlabel metal2 s 21270 29200 21326 30000 6 io_wbs_data_o[27]
port 25 nsew signal tristate
rlabel metal2 s 12254 0 12310 800 6 io_wbs_data_o[28]
port 26 nsew signal tristate
rlabel metal2 s 28354 29200 28410 30000 6 io_wbs_data_o[29]
port 27 nsew signal tristate
rlabel metal3 s 29200 27888 30000 28008 6 io_wbs_data_o[2]
port 28 nsew signal tristate
rlabel metal2 s 6458 0 6514 800 6 io_wbs_data_o[30]
port 29 nsew signal tristate
rlabel metal2 s 3238 0 3294 800 6 io_wbs_data_o[31]
port 30 nsew signal tristate
rlabel metal3 s 0 5448 800 5568 6 io_wbs_data_o[3]
port 31 nsew signal tristate
rlabel metal3 s 29200 29248 30000 29368 6 io_wbs_data_o[4]
port 32 nsew signal tristate
rlabel metal2 s 25134 29200 25190 30000 6 io_wbs_data_o[5]
port 33 nsew signal tristate
rlabel metal3 s 29200 688 30000 808 6 io_wbs_data_o[6]
port 34 nsew signal tristate
rlabel metal2 s 21914 0 21970 800 6 io_wbs_data_o[7]
port 35 nsew signal tristate
rlabel metal3 s 29200 12248 30000 12368 6 io_wbs_data_o[8]
port 36 nsew signal tristate
rlabel metal3 s 29200 8848 30000 8968 6 io_wbs_data_o[9]
port 37 nsew signal tristate
rlabel metal2 s 10322 29200 10378 30000 6 io_wbs_m2s_addr[0]
port 38 nsew signal input
rlabel metal2 s 11610 29200 11666 30000 6 io_wbs_m2s_addr[10]
port 39 nsew signal input
rlabel metal3 s 29200 21768 30000 21888 6 io_wbs_m2s_addr[11]
port 40 nsew signal input
rlabel metal3 s 0 4088 800 4208 6 io_wbs_m2s_addr[12]
port 41 nsew signal input
rlabel metal2 s 7746 0 7802 800 6 io_wbs_m2s_addr[13]
port 42 nsew signal input
rlabel metal3 s 29200 24488 30000 24608 6 io_wbs_m2s_addr[14]
port 43 nsew signal input
rlabel metal2 s 29642 0 29698 800 6 io_wbs_m2s_addr[15]
port 44 nsew signal input
rlabel metal2 s 17406 29200 17462 30000 6 io_wbs_m2s_addr[16]
port 45 nsew signal input
rlabel metal3 s 0 21768 800 21888 6 io_wbs_m2s_addr[17]
port 46 nsew signal input
rlabel metal2 s 8390 29200 8446 30000 6 io_wbs_m2s_addr[18]
port 47 nsew signal input
rlabel metal2 s 12898 29200 12954 30000 6 io_wbs_m2s_addr[19]
port 48 nsew signal input
rlabel metal3 s 29200 25168 30000 25288 6 io_wbs_m2s_addr[1]
port 49 nsew signal input
rlabel metal2 s 28998 0 29054 800 6 io_wbs_m2s_addr[20]
port 50 nsew signal input
rlabel metal2 s 14830 29200 14886 30000 6 io_wbs_m2s_addr[21]
port 51 nsew signal input
rlabel metal2 s 10966 0 11022 800 6 io_wbs_m2s_addr[22]
port 52 nsew signal input
rlabel metal3 s 29200 6808 30000 6928 6 io_wbs_m2s_addr[23]
port 53 nsew signal input
rlabel metal3 s 29200 18368 30000 18488 6 io_wbs_m2s_addr[24]
port 54 nsew signal input
rlabel metal3 s 0 14968 800 15088 6 io_wbs_m2s_addr[25]
port 55 nsew signal input
rlabel metal2 s 18050 29200 18106 30000 6 io_wbs_m2s_addr[26]
port 56 nsew signal input
rlabel metal2 s 5814 29200 5870 30000 6 io_wbs_m2s_addr[27]
port 57 nsew signal input
rlabel metal2 s 23202 0 23258 800 6 io_wbs_m2s_addr[28]
port 58 nsew signal input
rlabel metal3 s 0 3408 800 3528 6 io_wbs_m2s_addr[29]
port 59 nsew signal input
rlabel metal2 s 18694 0 18750 800 6 io_wbs_m2s_addr[2]
port 60 nsew signal input
rlabel metal2 s 1950 0 2006 800 6 io_wbs_m2s_addr[30]
port 61 nsew signal input
rlabel metal2 s 8390 0 8446 800 6 io_wbs_m2s_addr[31]
port 62 nsew signal input
rlabel metal2 s 27710 0 27766 800 6 io_wbs_m2s_addr[3]
port 63 nsew signal input
rlabel metal3 s 0 688 800 808 6 io_wbs_m2s_addr[4]
port 64 nsew signal input
rlabel metal3 s 29200 7488 30000 7608 6 io_wbs_m2s_addr[5]
port 65 nsew signal input
rlabel metal2 s 20626 0 20682 800 6 io_wbs_m2s_addr[6]
port 66 nsew signal input
rlabel metal3 s 0 24488 800 24608 6 io_wbs_m2s_addr[7]
port 67 nsew signal input
rlabel metal3 s 29200 2048 30000 2168 6 io_wbs_m2s_addr[8]
port 68 nsew signal input
rlabel metal3 s 0 6808 800 6928 6 io_wbs_m2s_addr[9]
port 69 nsew signal input
rlabel metal3 s 29200 11568 30000 11688 6 io_wbs_m2s_data[0]
port 70 nsew signal input
rlabel metal3 s 29200 19728 30000 19848 6 io_wbs_m2s_data[10]
port 71 nsew signal input
rlabel metal2 s 24490 0 24546 800 6 io_wbs_m2s_data[11]
port 72 nsew signal input
rlabel metal3 s 29200 21088 30000 21208 6 io_wbs_m2s_data[12]
port 73 nsew signal input
rlabel metal2 s 14186 0 14242 800 6 io_wbs_m2s_data[13]
port 74 nsew signal input
rlabel metal2 s 662 29200 718 30000 6 io_wbs_m2s_data[14]
port 75 nsew signal input
rlabel metal3 s 0 12928 800 13048 6 io_wbs_m2s_data[15]
port 76 nsew signal input
rlabel metal2 s 18 0 74 800 6 io_wbs_m2s_data[16]
port 77 nsew signal input
rlabel metal2 s 17406 0 17462 800 6 io_wbs_m2s_data[17]
port 78 nsew signal input
rlabel metal2 s 4526 29200 4582 30000 6 io_wbs_m2s_data[18]
port 79 nsew signal input
rlabel metal2 s 13542 29200 13598 30000 6 io_wbs_m2s_data[19]
port 80 nsew signal input
rlabel metal3 s 0 8168 800 8288 6 io_wbs_m2s_data[1]
port 81 nsew signal input
rlabel metal3 s 0 29248 800 29368 6 io_wbs_m2s_data[20]
port 82 nsew signal input
rlabel metal2 s 3882 0 3938 800 6 io_wbs_m2s_data[21]
port 83 nsew signal input
rlabel metal2 s 662 0 718 800 6 io_wbs_m2s_data[22]
port 84 nsew signal input
rlabel metal2 s 27066 29200 27122 30000 6 io_wbs_m2s_data[23]
port 85 nsew signal input
rlabel metal2 s 20626 29200 20682 30000 6 io_wbs_m2s_data[24]
port 86 nsew signal input
rlabel metal2 s 12898 0 12954 800 6 io_wbs_m2s_data[25]
port 87 nsew signal input
rlabel metal2 s 29642 29200 29698 30000 6 io_wbs_m2s_data[26]
port 88 nsew signal input
rlabel metal3 s 29200 3408 30000 3528 6 io_wbs_m2s_data[27]
port 89 nsew signal input
rlabel metal2 s 1306 29200 1362 30000 6 io_wbs_m2s_data[28]
port 90 nsew signal input
rlabel metal3 s 0 11568 800 11688 6 io_wbs_m2s_data[29]
port 91 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 io_wbs_m2s_data[2]
port 92 nsew signal input
rlabel metal2 s 9678 0 9734 800 6 io_wbs_m2s_data[30]
port 93 nsew signal input
rlabel metal2 s 15474 0 15530 800 6 io_wbs_m2s_data[31]
port 94 nsew signal input
rlabel metal3 s 29200 17008 30000 17128 6 io_wbs_m2s_data[3]
port 95 nsew signal input
rlabel metal2 s 16762 0 16818 800 6 io_wbs_m2s_data[4]
port 96 nsew signal input
rlabel metal2 s 23846 29200 23902 30000 6 io_wbs_m2s_data[5]
port 97 nsew signal input
rlabel metal2 s 22558 29200 22614 30000 6 io_wbs_m2s_data[6]
port 98 nsew signal input
rlabel metal2 s 2594 29200 2650 30000 6 io_wbs_m2s_data[7]
port 99 nsew signal input
rlabel metal2 s 7102 29200 7158 30000 6 io_wbs_m2s_data[8]
port 100 nsew signal input
rlabel metal2 s 19982 0 20038 800 6 io_wbs_m2s_data[9]
port 101 nsew signal input
rlabel metal3 s 0 8848 800 8968 6 io_wbs_m2s_stb
port 102 nsew signal input
rlabel metal3 s 0 26528 800 26648 6 io_wbs_m2s_we
port 103 nsew signal input
rlabel metal3 s 29200 13608 30000 13728 6 reset
port 104 nsew signal input
rlabel metal4 s 5576 2128 5896 27792 6 vccd1
port 105 nsew power input
rlabel metal4 s 14840 2128 15160 27792 6 vccd1
port 105 nsew power input
rlabel metal4 s 24104 2128 24424 27792 6 vccd1
port 105 nsew power input
rlabel metal4 s 10208 2128 10528 27792 6 vssd1
port 106 nsew ground input
rlabel metal4 s 19472 2128 19792 27792 6 vssd1
port 106 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 30000 30000
<< end >>
